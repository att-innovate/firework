// datapath.v

module datapath (
		input  wire [31:0] raw_data,
		input  wire        data_in_sel,
		input  wire        data_clr,
		input  wire        data_load,
		input  wire        data_out_sel,
		output wire        gt_eq_128,
		output wire [7:0]  encoded_byte
	);
	
	// TODO: implement datapath logic
	
endmodule
