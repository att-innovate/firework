// ghrd_10as066n2.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module ghrd_10as066n2 (
		input  wire        clk_100_clk,                                //                               clk_100.clk
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_ck,      //        emif_a10_hps_0_mem_conduit_end.mem_ck
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_ck_n,    //                                      .mem_ck_n
		output wire [16:0] emif_a10_hps_0_mem_conduit_end_mem_a,       //                                      .mem_a
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_act_n,   //                                      .mem_act_n
		output wire [1:0]  emif_a10_hps_0_mem_conduit_end_mem_ba,      //                                      .mem_ba
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_bg,      //                                      .mem_bg
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_cke,     //                                      .mem_cke
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_cs_n,    //                                      .mem_cs_n
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_odt,     //                                      .mem_odt
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_reset_n, //                                      .mem_reset_n
		output wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_par,     //                                      .mem_par
		input  wire [0:0]  emif_a10_hps_0_mem_conduit_end_mem_alert_n, //                                      .mem_alert_n
		inout  wire [3:0]  emif_a10_hps_0_mem_conduit_end_mem_dqs,     //                                      .mem_dqs
		inout  wire [3:0]  emif_a10_hps_0_mem_conduit_end_mem_dqs_n,   //                                      .mem_dqs_n
		inout  wire [31:0] emif_a10_hps_0_mem_conduit_end_mem_dq,      //                                      .mem_dq
		inout  wire [3:0]  emif_a10_hps_0_mem_conduit_end_mem_dbi_n,   //                                      .mem_dbi_n
		input  wire        emif_a10_hps_0_oct_conduit_end_oct_rzqin,   //        emif_a10_hps_0_oct_conduit_end.oct_rzqin
		input  wire        emif_a10_hps_0_pll_ref_clk_clock_sink_clk,  // emif_a10_hps_0_pll_ref_clk_clock_sink.clk
		input  wire        f2h_cold_reset_req_reset_n,                 //                    f2h_cold_reset_req.reset_n
		input  wire        f2h_debug_reset_req_reset_n,                //                   f2h_debug_reset_req.reset_n
		input  wire [27:0] f2h_stm_hw_events_stm_hwevents,             //                     f2h_stm_hw_events.stm_hwevents
		input  wire        f2h_warm_reset_req_reset_n,                 //                    f2h_warm_reset_req.reset_n
		output wire        hps_fpga_reset_reset,                       //                        hps_fpga_reset.reset
		output wire        hps_io_hps_io_phery_emac0_TX_CLK,           //                                hps_io.hps_io_phery_emac0_TX_CLK
		output wire        hps_io_hps_io_phery_emac0_TXD0,             //                                      .hps_io_phery_emac0_TXD0
		output wire        hps_io_hps_io_phery_emac0_TXD1,             //                                      .hps_io_phery_emac0_TXD1
		output wire        hps_io_hps_io_phery_emac0_TXD2,             //                                      .hps_io_phery_emac0_TXD2
		output wire        hps_io_hps_io_phery_emac0_TXD3,             //                                      .hps_io_phery_emac0_TXD3
		input  wire        hps_io_hps_io_phery_emac0_RX_CTL,           //                                      .hps_io_phery_emac0_RX_CTL
		output wire        hps_io_hps_io_phery_emac0_TX_CTL,           //                                      .hps_io_phery_emac0_TX_CTL
		input  wire        hps_io_hps_io_phery_emac0_RX_CLK,           //                                      .hps_io_phery_emac0_RX_CLK
		input  wire        hps_io_hps_io_phery_emac0_RXD0,             //                                      .hps_io_phery_emac0_RXD0
		input  wire        hps_io_hps_io_phery_emac0_RXD1,             //                                      .hps_io_phery_emac0_RXD1
		input  wire        hps_io_hps_io_phery_emac0_RXD2,             //                                      .hps_io_phery_emac0_RXD2
		input  wire        hps_io_hps_io_phery_emac0_RXD3,             //                                      .hps_io_phery_emac0_RXD3
		inout  wire        hps_io_hps_io_phery_emac0_MDIO,             //                                      .hps_io_phery_emac0_MDIO
		output wire        hps_io_hps_io_phery_emac0_MDC,              //                                      .hps_io_phery_emac0_MDC
		inout  wire        hps_io_hps_io_phery_sdmmc_CMD,              //                                      .hps_io_phery_sdmmc_CMD
		inout  wire        hps_io_hps_io_phery_sdmmc_D0,               //                                      .hps_io_phery_sdmmc_D0
		inout  wire        hps_io_hps_io_phery_sdmmc_D1,               //                                      .hps_io_phery_sdmmc_D1
		inout  wire        hps_io_hps_io_phery_sdmmc_D2,               //                                      .hps_io_phery_sdmmc_D2
		inout  wire        hps_io_hps_io_phery_sdmmc_D3,               //                                      .hps_io_phery_sdmmc_D3
		inout  wire        hps_io_hps_io_phery_sdmmc_D4,               //                                      .hps_io_phery_sdmmc_D4
		inout  wire        hps_io_hps_io_phery_sdmmc_D5,               //                                      .hps_io_phery_sdmmc_D5
		inout  wire        hps_io_hps_io_phery_sdmmc_D6,               //                                      .hps_io_phery_sdmmc_D6
		inout  wire        hps_io_hps_io_phery_sdmmc_D7,               //                                      .hps_io_phery_sdmmc_D7
		output wire        hps_io_hps_io_phery_sdmmc_CCLK,             //                                      .hps_io_phery_sdmmc_CCLK
		inout  wire        hps_io_hps_io_phery_usb0_DATA0,             //                                      .hps_io_phery_usb0_DATA0
		inout  wire        hps_io_hps_io_phery_usb0_DATA1,             //                                      .hps_io_phery_usb0_DATA1
		inout  wire        hps_io_hps_io_phery_usb0_DATA2,             //                                      .hps_io_phery_usb0_DATA2
		inout  wire        hps_io_hps_io_phery_usb0_DATA3,             //                                      .hps_io_phery_usb0_DATA3
		inout  wire        hps_io_hps_io_phery_usb0_DATA4,             //                                      .hps_io_phery_usb0_DATA4
		inout  wire        hps_io_hps_io_phery_usb0_DATA5,             //                                      .hps_io_phery_usb0_DATA5
		inout  wire        hps_io_hps_io_phery_usb0_DATA6,             //                                      .hps_io_phery_usb0_DATA6
		inout  wire        hps_io_hps_io_phery_usb0_DATA7,             //                                      .hps_io_phery_usb0_DATA7
		input  wire        hps_io_hps_io_phery_usb0_CLK,               //                                      .hps_io_phery_usb0_CLK
		output wire        hps_io_hps_io_phery_usb0_STP,               //                                      .hps_io_phery_usb0_STP
		input  wire        hps_io_hps_io_phery_usb0_DIR,               //                                      .hps_io_phery_usb0_DIR
		input  wire        hps_io_hps_io_phery_usb0_NXT,               //                                      .hps_io_phery_usb0_NXT
		output wire        hps_io_hps_io_phery_spim1_CLK,              //                                      .hps_io_phery_spim1_CLK
		output wire        hps_io_hps_io_phery_spim1_MOSI,             //                                      .hps_io_phery_spim1_MOSI
		input  wire        hps_io_hps_io_phery_spim1_MISO,             //                                      .hps_io_phery_spim1_MISO
		output wire        hps_io_hps_io_phery_spim1_SS0_N,            //                                      .hps_io_phery_spim1_SS0_N
		output wire        hps_io_hps_io_phery_spim1_SS1_N,            //                                      .hps_io_phery_spim1_SS1_N
		output wire        hps_io_hps_io_phery_trace_CLK,              //                                      .hps_io_phery_trace_CLK
		output wire        hps_io_hps_io_phery_trace_D0,               //                                      .hps_io_phery_trace_D0
		output wire        hps_io_hps_io_phery_trace_D1,               //                                      .hps_io_phery_trace_D1
		output wire        hps_io_hps_io_phery_trace_D2,               //                                      .hps_io_phery_trace_D2
		output wire        hps_io_hps_io_phery_trace_D3,               //                                      .hps_io_phery_trace_D3
		input  wire        hps_io_hps_io_phery_uart1_RX,               //                                      .hps_io_phery_uart1_RX
		output wire        hps_io_hps_io_phery_uart1_TX,               //                                      .hps_io_phery_uart1_TX
		inout  wire        hps_io_hps_io_phery_i2c1_SDA,               //                                      .hps_io_phery_i2c1_SDA
		inout  wire        hps_io_hps_io_phery_i2c1_SCL,               //                                      .hps_io_phery_i2c1_SCL
		inout  wire        hps_io_hps_io_gpio_gpio1_io5,               //                                      .hps_io_gpio_gpio1_io5
		inout  wire        hps_io_hps_io_gpio_gpio1_io14,              //                                      .hps_io_gpio_gpio1_io14
		inout  wire        hps_io_hps_io_gpio_gpio1_io16,              //                                      .hps_io_gpio_gpio1_io16
		inout  wire        hps_io_hps_io_gpio_gpio1_io17,              //                                      .hps_io_gpio_gpio1_io17
		output wire [2:0]  issp_hps_resets_source,                     //                       issp_hps_resets.source
		input  wire [3:0]  pio_button_external_connection_export,      //        pio_button_external_connection.export
		input  wire [3:0]  pio_dipsw_external_connection_export,       //         pio_dipsw_external_connection.export
		input  wire [3:0]  pio_led_external_connection_in_port,        //           pio_led_external_connection.in_port
		output wire [3:0]  pio_led_external_connection_out_port,       //                                      .out_port
		input  wire        reset_reset_n                               //                                 reset.reset_n
	);

	wire     [1:0] arria10_hps_0_emif_gp_to_emif;                         // arria10_hps_0:emif_gp_to_emif -> emif_a10_hps_0:hps_to_emif_gp
	wire  [4095:0] emif_a10_hps_0_hps_emif_conduit_end_emif_to_hps;       // emif_a10_hps_0:emif_to_hps -> arria10_hps_0:emif_emif_to_hps
	wire     [0:0] emif_a10_hps_0_hps_emif_conduit_end_emif_to_gp;        // emif_a10_hps_0:emif_to_hps_gp -> arria10_hps_0:emif_emif_to_gp
	wire  [4095:0] arria10_hps_0_emif_hps_to_emif;                        // arria10_hps_0:emif_hps_to_emif -> emif_a10_hps_0:hps_to_emif
	wire     [1:0] arria10_hps_0_h2f_axi_master_awburst;                  // arria10_hps_0:h2f_AWBURST -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awburst
	wire     [4:0] arria10_hps_0_h2f_axi_master_awuser;                   // arria10_hps_0:h2f_AWUSER -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awuser
	wire     [3:0] arria10_hps_0_h2f_axi_master_arlen;                    // arria10_hps_0:h2f_ARLEN -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arlen
	wire     [3:0] arria10_hps_0_h2f_axi_master_wstrb;                    // arria10_hps_0:h2f_WSTRB -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_wstrb
	wire           arria10_hps_0_h2f_axi_master_wready;                   // mm_interconnect_0:arria10_hps_0_h2f_axi_master_wready -> arria10_hps_0:h2f_WREADY
	wire     [3:0] arria10_hps_0_h2f_axi_master_rid;                      // mm_interconnect_0:arria10_hps_0_h2f_axi_master_rid -> arria10_hps_0:h2f_RID
	wire           arria10_hps_0_h2f_axi_master_rready;                   // arria10_hps_0:h2f_RREADY -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_rready
	wire     [3:0] arria10_hps_0_h2f_axi_master_awlen;                    // arria10_hps_0:h2f_AWLEN -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awlen
	wire     [3:0] arria10_hps_0_h2f_axi_master_wid;                      // arria10_hps_0:h2f_WID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_wid
	wire     [3:0] arria10_hps_0_h2f_axi_master_arcache;                  // arria10_hps_0:h2f_ARCACHE -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arcache
	wire           arria10_hps_0_h2f_axi_master_wvalid;                   // arria10_hps_0:h2f_WVALID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_wvalid
	wire    [31:0] arria10_hps_0_h2f_axi_master_araddr;                   // arria10_hps_0:h2f_ARADDR -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_araddr
	wire     [2:0] arria10_hps_0_h2f_axi_master_arprot;                   // arria10_hps_0:h2f_ARPROT -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arprot
	wire     [2:0] arria10_hps_0_h2f_axi_master_awprot;                   // arria10_hps_0:h2f_AWPROT -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awprot
	wire    [31:0] arria10_hps_0_h2f_axi_master_wdata;                    // arria10_hps_0:h2f_WDATA -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_wdata
	wire           arria10_hps_0_h2f_axi_master_arvalid;                  // arria10_hps_0:h2f_ARVALID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arvalid
	wire     [3:0] arria10_hps_0_h2f_axi_master_awcache;                  // arria10_hps_0:h2f_AWCACHE -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awcache
	wire     [3:0] arria10_hps_0_h2f_axi_master_arid;                     // arria10_hps_0:h2f_ARID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arid
	wire     [1:0] arria10_hps_0_h2f_axi_master_arlock;                   // arria10_hps_0:h2f_ARLOCK -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arlock
	wire     [1:0] arria10_hps_0_h2f_axi_master_awlock;                   // arria10_hps_0:h2f_AWLOCK -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awlock
	wire    [31:0] arria10_hps_0_h2f_axi_master_awaddr;                   // arria10_hps_0:h2f_AWADDR -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awaddr
	wire     [1:0] arria10_hps_0_h2f_axi_master_bresp;                    // mm_interconnect_0:arria10_hps_0_h2f_axi_master_bresp -> arria10_hps_0:h2f_BRESP
	wire           arria10_hps_0_h2f_axi_master_arready;                  // mm_interconnect_0:arria10_hps_0_h2f_axi_master_arready -> arria10_hps_0:h2f_ARREADY
	wire    [31:0] arria10_hps_0_h2f_axi_master_rdata;                    // mm_interconnect_0:arria10_hps_0_h2f_axi_master_rdata -> arria10_hps_0:h2f_RDATA
	wire           arria10_hps_0_h2f_axi_master_awready;                  // mm_interconnect_0:arria10_hps_0_h2f_axi_master_awready -> arria10_hps_0:h2f_AWREADY
	wire     [1:0] arria10_hps_0_h2f_axi_master_arburst;                  // arria10_hps_0:h2f_ARBURST -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arburst
	wire     [2:0] arria10_hps_0_h2f_axi_master_arsize;                   // arria10_hps_0:h2f_ARSIZE -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_arsize
	wire           arria10_hps_0_h2f_axi_master_bready;                   // arria10_hps_0:h2f_BREADY -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_bready
	wire           arria10_hps_0_h2f_axi_master_rlast;                    // mm_interconnect_0:arria10_hps_0_h2f_axi_master_rlast -> arria10_hps_0:h2f_RLAST
	wire           arria10_hps_0_h2f_axi_master_wlast;                    // arria10_hps_0:h2f_WLAST -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_wlast
	wire     [1:0] arria10_hps_0_h2f_axi_master_rresp;                    // mm_interconnect_0:arria10_hps_0_h2f_axi_master_rresp -> arria10_hps_0:h2f_RRESP
	wire     [3:0] arria10_hps_0_h2f_axi_master_awid;                     // arria10_hps_0:h2f_AWID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awid
	wire     [3:0] arria10_hps_0_h2f_axi_master_bid;                      // mm_interconnect_0:arria10_hps_0_h2f_axi_master_bid -> arria10_hps_0:h2f_BID
	wire           arria10_hps_0_h2f_axi_master_bvalid;                   // mm_interconnect_0:arria10_hps_0_h2f_axi_master_bvalid -> arria10_hps_0:h2f_BVALID
	wire     [2:0] arria10_hps_0_h2f_axi_master_awsize;                   // arria10_hps_0:h2f_AWSIZE -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awsize
	wire           arria10_hps_0_h2f_axi_master_awvalid;                  // arria10_hps_0:h2f_AWVALID -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_awvalid
	wire     [4:0] arria10_hps_0_h2f_axi_master_aruser;                   // arria10_hps_0:h2f_ARUSER -> mm_interconnect_0:arria10_hps_0_h2f_axi_master_aruser
	wire           arria10_hps_0_h2f_axi_master_rvalid;                   // mm_interconnect_0:arria10_hps_0_h2f_axi_master_rvalid -> arria10_hps_0:h2f_RVALID
	wire     [1:0] mm_interconnect_0_protobuf_serializer_0_s0_awburst;    // mm_interconnect_0:protobuf_serializer_0_s0_awburst -> protobuf_serializer_0:axs_s0_awburst
	wire     [7:0] mm_interconnect_0_protobuf_serializer_0_s0_arlen;      // mm_interconnect_0:protobuf_serializer_0_s0_arlen -> protobuf_serializer_0:axs_s0_arlen
	wire     [3:0] mm_interconnect_0_protobuf_serializer_0_s0_wstrb;      // mm_interconnect_0:protobuf_serializer_0_s0_wstrb -> protobuf_serializer_0:axs_s0_wstrb
	wire           mm_interconnect_0_protobuf_serializer_0_s0_wready;     // protobuf_serializer_0:axs_s0_wready -> mm_interconnect_0:protobuf_serializer_0_s0_wready
	wire     [3:0] mm_interconnect_0_protobuf_serializer_0_s0_rid;        // protobuf_serializer_0:axs_s0_rid -> mm_interconnect_0:protobuf_serializer_0_s0_rid
	wire           mm_interconnect_0_protobuf_serializer_0_s0_rready;     // mm_interconnect_0:protobuf_serializer_0_s0_rready -> protobuf_serializer_0:axs_s0_rready
	wire     [7:0] mm_interconnect_0_protobuf_serializer_0_s0_awlen;      // mm_interconnect_0:protobuf_serializer_0_s0_awlen -> protobuf_serializer_0:axs_s0_awlen
	wire           mm_interconnect_0_protobuf_serializer_0_s0_wvalid;     // mm_interconnect_0:protobuf_serializer_0_s0_wvalid -> protobuf_serializer_0:axs_s0_wvalid
	wire    [15:0] mm_interconnect_0_protobuf_serializer_0_s0_araddr;     // mm_interconnect_0:protobuf_serializer_0_s0_araddr -> protobuf_serializer_0:axs_s0_araddr
	wire    [31:0] mm_interconnect_0_protobuf_serializer_0_s0_wdata;      // mm_interconnect_0:protobuf_serializer_0_s0_wdata -> protobuf_serializer_0:axs_s0_wdata
	wire           mm_interconnect_0_protobuf_serializer_0_s0_arvalid;    // mm_interconnect_0:protobuf_serializer_0_s0_arvalid -> protobuf_serializer_0:axs_s0_arvalid
	wire     [3:0] mm_interconnect_0_protobuf_serializer_0_s0_arid;       // mm_interconnect_0:protobuf_serializer_0_s0_arid -> protobuf_serializer_0:axs_s0_arid
	wire    [15:0] mm_interconnect_0_protobuf_serializer_0_s0_awaddr;     // mm_interconnect_0:protobuf_serializer_0_s0_awaddr -> protobuf_serializer_0:axs_s0_awaddr
	wire           mm_interconnect_0_protobuf_serializer_0_s0_arready;    // protobuf_serializer_0:axs_s0_arready -> mm_interconnect_0:protobuf_serializer_0_s0_arready
	wire    [31:0] mm_interconnect_0_protobuf_serializer_0_s0_rdata;      // protobuf_serializer_0:axs_s0_rdata -> mm_interconnect_0:protobuf_serializer_0_s0_rdata
	wire           mm_interconnect_0_protobuf_serializer_0_s0_awready;    // protobuf_serializer_0:axs_s0_awready -> mm_interconnect_0:protobuf_serializer_0_s0_awready
	wire     [1:0] mm_interconnect_0_protobuf_serializer_0_s0_arburst;    // mm_interconnect_0:protobuf_serializer_0_s0_arburst -> protobuf_serializer_0:axs_s0_arburst
	wire     [2:0] mm_interconnect_0_protobuf_serializer_0_s0_arsize;     // mm_interconnect_0:protobuf_serializer_0_s0_arsize -> protobuf_serializer_0:axs_s0_arsize
	wire           mm_interconnect_0_protobuf_serializer_0_s0_bready;     // mm_interconnect_0:protobuf_serializer_0_s0_bready -> protobuf_serializer_0:axs_s0_bready
	wire           mm_interconnect_0_protobuf_serializer_0_s0_rlast;      // protobuf_serializer_0:axs_s0_rlast -> mm_interconnect_0:protobuf_serializer_0_s0_rlast
	wire     [3:0] mm_interconnect_0_protobuf_serializer_0_s0_awid;       // mm_interconnect_0:protobuf_serializer_0_s0_awid -> protobuf_serializer_0:axs_s0_awid
	wire     [3:0] mm_interconnect_0_protobuf_serializer_0_s0_bid;        // protobuf_serializer_0:axs_s0_bid -> mm_interconnect_0:protobuf_serializer_0_s0_bid
	wire           mm_interconnect_0_protobuf_serializer_0_s0_bvalid;     // protobuf_serializer_0:axs_s0_bvalid -> mm_interconnect_0:protobuf_serializer_0_s0_bvalid
	wire     [2:0] mm_interconnect_0_protobuf_serializer_0_s0_awsize;     // mm_interconnect_0:protobuf_serializer_0_s0_awsize -> protobuf_serializer_0:axs_s0_awsize
	wire           mm_interconnect_0_protobuf_serializer_0_s0_awvalid;    // mm_interconnect_0:protobuf_serializer_0_s0_awvalid -> protobuf_serializer_0:axs_s0_awvalid
	wire           mm_interconnect_0_protobuf_serializer_0_s0_rvalid;     // protobuf_serializer_0:axs_s0_rvalid -> mm_interconnect_0:protobuf_serializer_0_s0_rvalid
	wire           mm_interconnect_0_onchip_memory2_0_s1_chipselect;      // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire     [7:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;        // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire    [17:0] mm_interconnect_0_onchip_memory2_0_s1_address;         // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire           mm_interconnect_0_onchip_memory2_0_s1_write;           // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire     [7:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;       // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire           mm_interconnect_0_onchip_memory2_0_s1_clken;           // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_awburst;               // arria10_hps_0:h2f_lw_AWBURST -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awburst
	wire     [4:0] arria10_hps_0_h2f_lw_axi_master_awuser;                // arria10_hps_0:h2f_lw_AWUSER -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awuser
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_arlen;                 // arria10_hps_0:h2f_lw_ARLEN -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arlen
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_wstrb;                 // arria10_hps_0:h2f_lw_WSTRB -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wstrb
	wire           arria10_hps_0_h2f_lw_axi_master_wready;                // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wready -> arria10_hps_0:h2f_lw_WREADY
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_rid;                   // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rid -> arria10_hps_0:h2f_lw_RID
	wire           arria10_hps_0_h2f_lw_axi_master_rready;                // arria10_hps_0:h2f_lw_RREADY -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rready
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_awlen;                 // arria10_hps_0:h2f_lw_AWLEN -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awlen
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_wid;                   // arria10_hps_0:h2f_lw_WID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wid
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_arcache;               // arria10_hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arcache
	wire           arria10_hps_0_h2f_lw_axi_master_wvalid;                // arria10_hps_0:h2f_lw_WVALID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wvalid
	wire    [20:0] arria10_hps_0_h2f_lw_axi_master_araddr;                // arria10_hps_0:h2f_lw_ARADDR -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_araddr
	wire     [2:0] arria10_hps_0_h2f_lw_axi_master_arprot;                // arria10_hps_0:h2f_lw_ARPROT -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arprot
	wire     [2:0] arria10_hps_0_h2f_lw_axi_master_awprot;                // arria10_hps_0:h2f_lw_AWPROT -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awprot
	wire    [31:0] arria10_hps_0_h2f_lw_axi_master_wdata;                 // arria10_hps_0:h2f_lw_WDATA -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wdata
	wire           arria10_hps_0_h2f_lw_axi_master_arvalid;               // arria10_hps_0:h2f_lw_ARVALID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arvalid
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_awcache;               // arria10_hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awcache
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_arid;                  // arria10_hps_0:h2f_lw_ARID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arid
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_arlock;                // arria10_hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arlock
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_awlock;                // arria10_hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awlock
	wire    [20:0] arria10_hps_0_h2f_lw_axi_master_awaddr;                // arria10_hps_0:h2f_lw_AWADDR -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awaddr
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_bresp;                 // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_bresp -> arria10_hps_0:h2f_lw_BRESP
	wire           arria10_hps_0_h2f_lw_axi_master_arready;               // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arready -> arria10_hps_0:h2f_lw_ARREADY
	wire    [31:0] arria10_hps_0_h2f_lw_axi_master_rdata;                 // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rdata -> arria10_hps_0:h2f_lw_RDATA
	wire           arria10_hps_0_h2f_lw_axi_master_awready;               // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awready -> arria10_hps_0:h2f_lw_AWREADY
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_arburst;               // arria10_hps_0:h2f_lw_ARBURST -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arburst
	wire     [2:0] arria10_hps_0_h2f_lw_axi_master_arsize;                // arria10_hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_arsize
	wire           arria10_hps_0_h2f_lw_axi_master_bready;                // arria10_hps_0:h2f_lw_BREADY -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_bready
	wire           arria10_hps_0_h2f_lw_axi_master_rlast;                 // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rlast -> arria10_hps_0:h2f_lw_RLAST
	wire           arria10_hps_0_h2f_lw_axi_master_wlast;                 // arria10_hps_0:h2f_lw_WLAST -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_wlast
	wire     [1:0] arria10_hps_0_h2f_lw_axi_master_rresp;                 // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rresp -> arria10_hps_0:h2f_lw_RRESP
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_awid;                  // arria10_hps_0:h2f_lw_AWID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awid
	wire     [3:0] arria10_hps_0_h2f_lw_axi_master_bid;                   // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_bid -> arria10_hps_0:h2f_lw_BID
	wire           arria10_hps_0_h2f_lw_axi_master_bvalid;                // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_bvalid -> arria10_hps_0:h2f_lw_BVALID
	wire     [2:0] arria10_hps_0_h2f_lw_axi_master_awsize;                // arria10_hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awsize
	wire           arria10_hps_0_h2f_lw_axi_master_awvalid;               // arria10_hps_0:h2f_lw_AWVALID -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_awvalid
	wire     [4:0] arria10_hps_0_h2f_lw_axi_master_aruser;                // arria10_hps_0:h2f_lw_ARUSER -> mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_aruser
	wire           arria10_hps_0_h2f_lw_axi_master_rvalid;                // mm_interconnect_1:arria10_hps_0_h2f_lw_axi_master_rvalid -> arria10_hps_0:h2f_lw_RVALID
	wire    [31:0] fpga_only_master_master_readdata;                      // mm_interconnect_1:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire           fpga_only_master_master_waitrequest;                   // mm_interconnect_1:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire    [31:0] fpga_only_master_master_address;                       // fpga_only_master:master_address -> mm_interconnect_1:fpga_only_master_master_address
	wire           fpga_only_master_master_read;                          // fpga_only_master:master_read -> mm_interconnect_1:fpga_only_master_master_read
	wire     [3:0] fpga_only_master_master_byteenable;                    // fpga_only_master:master_byteenable -> mm_interconnect_1:fpga_only_master_master_byteenable
	wire           fpga_only_master_master_readdatavalid;                 // mm_interconnect_1:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire           fpga_only_master_master_write;                         // fpga_only_master:master_write -> mm_interconnect_1:fpga_only_master_master_write
	wire    [31:0] fpga_only_master_master_writedata;                     // fpga_only_master:master_writedata -> mm_interconnect_1:fpga_only_master_master_writedata
	wire    [31:0] mm_interconnect_1_pb_lwh2f_s0_readdata;                // pb_lwh2f:s0_readdata -> mm_interconnect_1:pb_lwh2f_s0_readdata
	wire           mm_interconnect_1_pb_lwh2f_s0_waitrequest;             // pb_lwh2f:s0_waitrequest -> mm_interconnect_1:pb_lwh2f_s0_waitrequest
	wire           mm_interconnect_1_pb_lwh2f_s0_debugaccess;             // mm_interconnect_1:pb_lwh2f_s0_debugaccess -> pb_lwh2f:s0_debugaccess
	wire     [8:0] mm_interconnect_1_pb_lwh2f_s0_address;                 // mm_interconnect_1:pb_lwh2f_s0_address -> pb_lwh2f:s0_address
	wire           mm_interconnect_1_pb_lwh2f_s0_read;                    // mm_interconnect_1:pb_lwh2f_s0_read -> pb_lwh2f:s0_read
	wire     [3:0] mm_interconnect_1_pb_lwh2f_s0_byteenable;              // mm_interconnect_1:pb_lwh2f_s0_byteenable -> pb_lwh2f:s0_byteenable
	wire           mm_interconnect_1_pb_lwh2f_s0_readdatavalid;           // pb_lwh2f:s0_readdatavalid -> mm_interconnect_1:pb_lwh2f_s0_readdatavalid
	wire           mm_interconnect_1_pb_lwh2f_s0_write;                   // mm_interconnect_1:pb_lwh2f_s0_write -> pb_lwh2f:s0_write
	wire    [31:0] mm_interconnect_1_pb_lwh2f_s0_writedata;               // mm_interconnect_1:pb_lwh2f_s0_writedata -> pb_lwh2f:s0_writedata
	wire     [0:0] mm_interconnect_1_pb_lwh2f_s0_burstcount;              // mm_interconnect_1:pb_lwh2f_s0_burstcount -> pb_lwh2f:s0_burstcount
	wire           pb_lwh2f_m0_waitrequest;                               // mm_interconnect_2:pb_lwh2f_m0_waitrequest -> pb_lwh2f:m0_waitrequest
	wire    [31:0] pb_lwh2f_m0_readdata;                                  // mm_interconnect_2:pb_lwh2f_m0_readdata -> pb_lwh2f:m0_readdata
	wire           pb_lwh2f_m0_debugaccess;                               // pb_lwh2f:m0_debugaccess -> mm_interconnect_2:pb_lwh2f_m0_debugaccess
	wire     [8:0] pb_lwh2f_m0_address;                                   // pb_lwh2f:m0_address -> mm_interconnect_2:pb_lwh2f_m0_address
	wire           pb_lwh2f_m0_read;                                      // pb_lwh2f:m0_read -> mm_interconnect_2:pb_lwh2f_m0_read
	wire     [3:0] pb_lwh2f_m0_byteenable;                                // pb_lwh2f:m0_byteenable -> mm_interconnect_2:pb_lwh2f_m0_byteenable
	wire           pb_lwh2f_m0_readdatavalid;                             // mm_interconnect_2:pb_lwh2f_m0_readdatavalid -> pb_lwh2f:m0_readdatavalid
	wire    [31:0] pb_lwh2f_m0_writedata;                                 // pb_lwh2f:m0_writedata -> mm_interconnect_2:pb_lwh2f_m0_writedata
	wire           pb_lwh2f_m0_write;                                     // pb_lwh2f:m0_write -> mm_interconnect_2:pb_lwh2f_m0_write
	wire     [0:0] pb_lwh2f_m0_burstcount;                                // pb_lwh2f:m0_burstcount -> mm_interconnect_2:pb_lwh2f_m0_burstcount
	wire    [31:0] mm_interconnect_2_ilc_avalon_slave_readdata;           // ILC:avmm_rddata -> mm_interconnect_2:ILC_avalon_slave_readdata
	wire     [5:0] mm_interconnect_2_ilc_avalon_slave_address;            // mm_interconnect_2:ILC_avalon_slave_address -> ILC:avmm_addr
	wire           mm_interconnect_2_ilc_avalon_slave_read;               // mm_interconnect_2:ILC_avalon_slave_read -> ILC:avmm_read
	wire           mm_interconnect_2_ilc_avalon_slave_write;              // mm_interconnect_2:ILC_avalon_slave_write -> ILC:avmm_write
	wire    [31:0] mm_interconnect_2_ilc_avalon_slave_writedata;          // mm_interconnect_2:ILC_avalon_slave_writedata -> ILC:avmm_wrdata
	wire    [31:0] mm_interconnect_2_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_2:sysid_qsys_0_control_slave_readdata
	wire     [0:0] mm_interconnect_2_sysid_qsys_0_control_slave_address;  // mm_interconnect_2:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire           mm_interconnect_2_led_pio_s1_chipselect;               // mm_interconnect_2:led_pio_s1_chipselect -> led_pio:chipselect
	wire    [31:0] mm_interconnect_2_led_pio_s1_readdata;                 // led_pio:readdata -> mm_interconnect_2:led_pio_s1_readdata
	wire     [1:0] mm_interconnect_2_led_pio_s1_address;                  // mm_interconnect_2:led_pio_s1_address -> led_pio:address
	wire           mm_interconnect_2_led_pio_s1_write;                    // mm_interconnect_2:led_pio_s1_write -> led_pio:write_n
	wire    [31:0] mm_interconnect_2_led_pio_s1_writedata;                // mm_interconnect_2:led_pio_s1_writedata -> led_pio:writedata
	wire           mm_interconnect_2_button_pio_s1_chipselect;            // mm_interconnect_2:button_pio_s1_chipselect -> button_pio:chipselect
	wire    [31:0] mm_interconnect_2_button_pio_s1_readdata;              // button_pio:readdata -> mm_interconnect_2:button_pio_s1_readdata
	wire     [1:0] mm_interconnect_2_button_pio_s1_address;               // mm_interconnect_2:button_pio_s1_address -> button_pio:address
	wire           mm_interconnect_2_button_pio_s1_write;                 // mm_interconnect_2:button_pio_s1_write -> button_pio:write_n
	wire    [31:0] mm_interconnect_2_button_pio_s1_writedata;             // mm_interconnect_2:button_pio_s1_writedata -> button_pio:writedata
	wire           mm_interconnect_2_dipsw_pio_s1_chipselect;             // mm_interconnect_2:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire    [31:0] mm_interconnect_2_dipsw_pio_s1_readdata;               // dipsw_pio:readdata -> mm_interconnect_2:dipsw_pio_s1_readdata
	wire     [1:0] mm_interconnect_2_dipsw_pio_s1_address;                // mm_interconnect_2:dipsw_pio_s1_address -> dipsw_pio:address
	wire           mm_interconnect_2_dipsw_pio_s1_write;                  // mm_interconnect_2:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire    [31:0] mm_interconnect_2_dipsw_pio_s1_writedata;              // mm_interconnect_2:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire    [31:0] hps_only_master_master_readdata;                       // mm_interconnect_3:hps_only_master_master_readdata -> hps_only_master:master_readdata
	wire           hps_only_master_master_waitrequest;                    // mm_interconnect_3:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	wire    [31:0] hps_only_master_master_address;                        // hps_only_master:master_address -> mm_interconnect_3:hps_only_master_master_address
	wire           hps_only_master_master_read;                           // hps_only_master:master_read -> mm_interconnect_3:hps_only_master_master_read
	wire     [3:0] hps_only_master_master_byteenable;                     // hps_only_master:master_byteenable -> mm_interconnect_3:hps_only_master_master_byteenable
	wire           hps_only_master_master_readdatavalid;                  // mm_interconnect_3:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	wire           hps_only_master_master_write;                          // hps_only_master:master_write -> mm_interconnect_3:hps_only_master_master_write
	wire    [31:0] hps_only_master_master_writedata;                      // hps_only_master:master_writedata -> mm_interconnect_3:hps_only_master_master_writedata
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awburst; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awburst -> arria10_hps_0:f2h_AWBURST
	wire     [4:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awuser;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awuser -> arria10_hps_0:f2h_AWUSER
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlen;   // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arlen -> arria10_hps_0:f2h_ARLEN
	wire    [15:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wstrb;   // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wstrb -> arria10_hps_0:f2h_WSTRB
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wready;  // arria10_hps_0:f2h_WREADY -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wready
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rid;     // arria10_hps_0:f2h_RID -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rid
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rready;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rready -> arria10_hps_0:f2h_RREADY
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlen;   // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awlen -> arria10_hps_0:f2h_AWLEN
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wid;     // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wid -> arria10_hps_0:f2h_WID
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arcache; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arcache -> arria10_hps_0:f2h_ARCACHE
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wvalid;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wvalid -> arria10_hps_0:f2h_WVALID
	wire    [31:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_araddr;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_araddr -> arria10_hps_0:f2h_ARADDR
	wire     [2:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arprot;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arprot -> arria10_hps_0:f2h_ARPROT
	wire     [2:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awprot;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awprot -> arria10_hps_0:f2h_AWPROT
	wire   [127:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wdata;   // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wdata -> arria10_hps_0:f2h_WDATA
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arvalid; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arvalid -> arria10_hps_0:f2h_ARVALID
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awcache; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awcache -> arria10_hps_0:f2h_AWCACHE
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arid;    // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arid -> arria10_hps_0:f2h_ARID
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlock;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arlock -> arria10_hps_0:f2h_ARLOCK
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlock;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awlock -> arria10_hps_0:f2h_AWLOCK
	wire    [31:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awaddr;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awaddr -> arria10_hps_0:f2h_AWADDR
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bresp;   // arria10_hps_0:f2h_BRESP -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_bresp
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arready; // arria10_hps_0:f2h_ARREADY -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arready
	wire   [127:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rdata;   // arria10_hps_0:f2h_RDATA -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rdata
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awready; // arria10_hps_0:f2h_AWREADY -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awready
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arburst; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arburst -> arria10_hps_0:f2h_ARBURST
	wire     [2:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arsize;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_arsize -> arria10_hps_0:f2h_ARSIZE
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bready;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_bready -> arria10_hps_0:f2h_BREADY
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rlast;   // arria10_hps_0:f2h_RLAST -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rlast
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wlast;   // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_wlast -> arria10_hps_0:f2h_WLAST
	wire     [1:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rresp;   // arria10_hps_0:f2h_RRESP -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rresp
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awid;    // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awid -> arria10_hps_0:f2h_AWID
	wire     [3:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bid;     // arria10_hps_0:f2h_BID -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_bid
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bvalid;  // arria10_hps_0:f2h_BVALID -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_bvalid
	wire     [2:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awsize;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awsize -> arria10_hps_0:f2h_AWSIZE
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awvalid; // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_awvalid -> arria10_hps_0:f2h_AWVALID
	wire     [4:0] mm_interconnect_3_arria10_hps_0_f2h_axi_slave_aruser;  // mm_interconnect_3:arria10_hps_0_f2h_axi_slave_aruser -> arria10_hps_0:f2h_ARUSER
	wire           mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rvalid;  // arria10_hps_0:f2h_RVALID -> mm_interconnect_3:arria10_hps_0_f2h_axi_slave_rvalid
	wire    [31:0] f2sdram_only_master1_master_readdata;                  // mm_interconnect_4:f2sdram_only_master1_master_readdata -> f2sdram_only_master1:master_readdata
	wire           f2sdram_only_master1_master_waitrequest;               // mm_interconnect_4:f2sdram_only_master1_master_waitrequest -> f2sdram_only_master1:master_waitrequest
	wire    [31:0] f2sdram_only_master1_master_address;                   // f2sdram_only_master1:master_address -> mm_interconnect_4:f2sdram_only_master1_master_address
	wire           f2sdram_only_master1_master_read;                      // f2sdram_only_master1:master_read -> mm_interconnect_4:f2sdram_only_master1_master_read
	wire     [3:0] f2sdram_only_master1_master_byteenable;                // f2sdram_only_master1:master_byteenable -> mm_interconnect_4:f2sdram_only_master1_master_byteenable
	wire           f2sdram_only_master1_master_readdatavalid;             // mm_interconnect_4:f2sdram_only_master1_master_readdatavalid -> f2sdram_only_master1:master_readdatavalid
	wire           f2sdram_only_master1_master_write;                     // f2sdram_only_master1:master_write -> mm_interconnect_4:f2sdram_only_master1_master_write
	wire    [31:0] f2sdram_only_master1_master_writedata;                 // f2sdram_only_master1:master_writedata -> mm_interconnect_4:f2sdram_only_master1_master_writedata
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awburst; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awburst -> arria10_hps_0:f2sdram0_AWBURST
	wire     [4:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awuser;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awuser -> arria10_hps_0:f2sdram0_AWUSER
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlen;   // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arlen -> arria10_hps_0:f2sdram0_ARLEN
	wire    [15:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_wstrb;   // mm_interconnect_4:arria10_hps_0_f2sdram0_data_wstrb -> arria10_hps_0:f2sdram0_WSTRB
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_wready;  // arria10_hps_0:f2sdram0_WREADY -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_wready
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_rid;     // arria10_hps_0:f2sdram0_RID -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_rid
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_rready;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_rready -> arria10_hps_0:f2sdram0_RREADY
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlen;   // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awlen -> arria10_hps_0:f2sdram0_AWLEN
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_wid;     // mm_interconnect_4:arria10_hps_0_f2sdram0_data_wid -> arria10_hps_0:f2sdram0_WID
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arcache; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arcache -> arria10_hps_0:f2sdram0_ARCACHE
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_wvalid;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_wvalid -> arria10_hps_0:f2sdram0_WVALID
	wire    [31:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_araddr;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_araddr -> arria10_hps_0:f2sdram0_ARADDR
	wire     [2:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arprot;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arprot -> arria10_hps_0:f2sdram0_ARPROT
	wire     [2:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awprot;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awprot -> arria10_hps_0:f2sdram0_AWPROT
	wire   [127:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_wdata;   // mm_interconnect_4:arria10_hps_0_f2sdram0_data_wdata -> arria10_hps_0:f2sdram0_WDATA
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_arvalid; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arvalid -> arria10_hps_0:f2sdram0_ARVALID
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awcache; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awcache -> arria10_hps_0:f2sdram0_AWCACHE
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arid;    // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arid -> arria10_hps_0:f2sdram0_ARID
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlock;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arlock -> arria10_hps_0:f2sdram0_ARLOCK
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlock;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awlock -> arria10_hps_0:f2sdram0_AWLOCK
	wire    [31:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awaddr;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awaddr -> arria10_hps_0:f2sdram0_AWADDR
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_bresp;   // arria10_hps_0:f2sdram0_BRESP -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_bresp
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_arready; // arria10_hps_0:f2sdram0_ARREADY -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_arready
	wire   [127:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_rdata;   // arria10_hps_0:f2sdram0_RDATA -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_rdata
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_awready; // arria10_hps_0:f2sdram0_AWREADY -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_awready
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arburst; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arburst -> arria10_hps_0:f2sdram0_ARBURST
	wire     [2:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_arsize;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_arsize -> arria10_hps_0:f2sdram0_ARSIZE
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_bready;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_bready -> arria10_hps_0:f2sdram0_BREADY
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_rlast;   // arria10_hps_0:f2sdram0_RLAST -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_rlast
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_wlast;   // mm_interconnect_4:arria10_hps_0_f2sdram0_data_wlast -> arria10_hps_0:f2sdram0_WLAST
	wire     [1:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_rresp;   // arria10_hps_0:f2sdram0_RRESP -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_rresp
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awid;    // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awid -> arria10_hps_0:f2sdram0_AWID
	wire     [3:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_bid;     // arria10_hps_0:f2sdram0_BID -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_bid
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_bvalid;  // arria10_hps_0:f2sdram0_BVALID -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_bvalid
	wire     [2:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_awsize;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awsize -> arria10_hps_0:f2sdram0_AWSIZE
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_awvalid; // mm_interconnect_4:arria10_hps_0_f2sdram0_data_awvalid -> arria10_hps_0:f2sdram0_AWVALID
	wire     [4:0] mm_interconnect_4_arria10_hps_0_f2sdram0_data_aruser;  // mm_interconnect_4:arria10_hps_0_f2sdram0_data_aruser -> arria10_hps_0:f2sdram0_ARUSER
	wire           mm_interconnect_4_arria10_hps_0_f2sdram0_data_rvalid;  // arria10_hps_0:f2sdram0_RVALID -> mm_interconnect_4:arria10_hps_0_f2sdram0_data_rvalid
	wire    [31:0] f2sdram_only_master_master_readdata;                   // mm_interconnect_5:f2sdram_only_master_master_readdata -> f2sdram_only_master:master_readdata
	wire           f2sdram_only_master_master_waitrequest;                // mm_interconnect_5:f2sdram_only_master_master_waitrequest -> f2sdram_only_master:master_waitrequest
	wire    [31:0] f2sdram_only_master_master_address;                    // f2sdram_only_master:master_address -> mm_interconnect_5:f2sdram_only_master_master_address
	wire           f2sdram_only_master_master_read;                       // f2sdram_only_master:master_read -> mm_interconnect_5:f2sdram_only_master_master_read
	wire     [3:0] f2sdram_only_master_master_byteenable;                 // f2sdram_only_master:master_byteenable -> mm_interconnect_5:f2sdram_only_master_master_byteenable
	wire           f2sdram_only_master_master_readdatavalid;              // mm_interconnect_5:f2sdram_only_master_master_readdatavalid -> f2sdram_only_master:master_readdatavalid
	wire           f2sdram_only_master_master_write;                      // f2sdram_only_master:master_write -> mm_interconnect_5:f2sdram_only_master_master_write
	wire    [31:0] f2sdram_only_master_master_writedata;                  // f2sdram_only_master:master_writedata -> mm_interconnect_5:f2sdram_only_master_master_writedata
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awburst; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awburst -> arria10_hps_0:f2sdram2_AWBURST
	wire     [4:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awuser;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awuser -> arria10_hps_0:f2sdram2_AWUSER
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlen;   // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arlen -> arria10_hps_0:f2sdram2_ARLEN
	wire    [15:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_wstrb;   // mm_interconnect_5:arria10_hps_0_f2sdram2_data_wstrb -> arria10_hps_0:f2sdram2_WSTRB
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_wready;  // arria10_hps_0:f2sdram2_WREADY -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_wready
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_rid;     // arria10_hps_0:f2sdram2_RID -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_rid
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_rready;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_rready -> arria10_hps_0:f2sdram2_RREADY
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlen;   // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awlen -> arria10_hps_0:f2sdram2_AWLEN
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_wid;     // mm_interconnect_5:arria10_hps_0_f2sdram2_data_wid -> arria10_hps_0:f2sdram2_WID
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arcache; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arcache -> arria10_hps_0:f2sdram2_ARCACHE
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_wvalid;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_wvalid -> arria10_hps_0:f2sdram2_WVALID
	wire    [31:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_araddr;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_araddr -> arria10_hps_0:f2sdram2_ARADDR
	wire     [2:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arprot;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arprot -> arria10_hps_0:f2sdram2_ARPROT
	wire     [2:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awprot;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awprot -> arria10_hps_0:f2sdram2_AWPROT
	wire   [127:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_wdata;   // mm_interconnect_5:arria10_hps_0_f2sdram2_data_wdata -> arria10_hps_0:f2sdram2_WDATA
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_arvalid; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arvalid -> arria10_hps_0:f2sdram2_ARVALID
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awcache; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awcache -> arria10_hps_0:f2sdram2_AWCACHE
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arid;    // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arid -> arria10_hps_0:f2sdram2_ARID
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlock;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arlock -> arria10_hps_0:f2sdram2_ARLOCK
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlock;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awlock -> arria10_hps_0:f2sdram2_AWLOCK
	wire    [31:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awaddr;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awaddr -> arria10_hps_0:f2sdram2_AWADDR
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_bresp;   // arria10_hps_0:f2sdram2_BRESP -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_bresp
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_arready; // arria10_hps_0:f2sdram2_ARREADY -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_arready
	wire   [127:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_rdata;   // arria10_hps_0:f2sdram2_RDATA -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_rdata
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_awready; // arria10_hps_0:f2sdram2_AWREADY -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_awready
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arburst; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arburst -> arria10_hps_0:f2sdram2_ARBURST
	wire     [2:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_arsize;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_arsize -> arria10_hps_0:f2sdram2_ARSIZE
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_bready;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_bready -> arria10_hps_0:f2sdram2_BREADY
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_rlast;   // arria10_hps_0:f2sdram2_RLAST -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_rlast
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_wlast;   // mm_interconnect_5:arria10_hps_0_f2sdram2_data_wlast -> arria10_hps_0:f2sdram2_WLAST
	wire     [1:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_rresp;   // arria10_hps_0:f2sdram2_RRESP -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_rresp
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awid;    // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awid -> arria10_hps_0:f2sdram2_AWID
	wire     [3:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_bid;     // arria10_hps_0:f2sdram2_BID -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_bid
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_bvalid;  // arria10_hps_0:f2sdram2_BVALID -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_bvalid
	wire     [2:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_awsize;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awsize -> arria10_hps_0:f2sdram2_AWSIZE
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_awvalid; // mm_interconnect_5:arria10_hps_0_f2sdram2_data_awvalid -> arria10_hps_0:f2sdram2_AWVALID
	wire     [4:0] mm_interconnect_5_arria10_hps_0_f2sdram2_data_aruser;  // mm_interconnect_5:arria10_hps_0_f2sdram2_data_aruser -> arria10_hps_0:f2sdram2_ARUSER
	wire           mm_interconnect_5_arria10_hps_0_f2sdram2_data_rvalid;  // arria10_hps_0:f2sdram2_RVALID -> mm_interconnect_5:arria10_hps_0_f2sdram2_data_rvalid
	wire     [1:0] ilc_irq_irq;                                           // irq_mapper:sender_irq -> ILC:irq
	wire    [31:0] arria10_hps_0_f2h_irq0_irq;                            // irq_mapper_001:sender_irq -> arria10_hps_0:f2h_irq_p0
	wire    [31:0] arria10_hps_0_f2h_irq1_irq;                            // irq_mapper_002:sender_irq -> arria10_hps_0:f2h_irq_p1
	wire           irq_mapper_receiver0_irq;                              // button_pio:irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire           irq_mapper_receiver1_irq;                              // dipsw_pio:irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire           rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire           arria10_hps_0_h2f_reset_reset;                         // arria10_hps_0:h2f_rst_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1]
	wire           rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> f2sdram_only_master:clk_reset_reset
	wire           rst_controller_002_reset_out_reset;                    // rst_controller_002:reset_out -> f2sdram_only_master1:clk_reset_reset
	wire           rst_controller_003_reset_out_reset;                    // rst_controller_003:reset_out -> fpga_only_master:clk_reset_reset
	wire           rst_controller_004_reset_out_reset;                    // rst_controller_004:reset_out -> hps_only_master:clk_reset_reset

	interrupt_latency_counter #(
		.INTR_TYPE    (0),
		.CLOCK_RATE   (100000000),
		.IRQ_PORT_CNT (2)
	) ilc (
		.reset_n     (~hps_fpga_reset_reset),                        //      reset_n.reset_n
		.clk         (clk_100_clk),                                  //          clk.clk
		.irq         (ilc_irq_irq),                                  //          irq.irq
		.avmm_addr   (mm_interconnect_2_ilc_avalon_slave_address),   // avalon_slave.address
		.avmm_wrdata (mm_interconnect_2_ilc_avalon_slave_writedata), //             .writedata
		.avmm_write  (mm_interconnect_2_ilc_avalon_slave_write),     //             .write
		.avmm_read   (mm_interconnect_2_ilc_avalon_slave_read),      //             .read
		.avmm_rddata (mm_interconnect_2_ilc_avalon_slave_readdata)   //             .readdata
	);

	ghrd_10as066n2_altera_arria10_hps_161_wdommvq #(
		.F2S_Width (6),
		.S2F_Width (4)
	) arria10_hps_0 (
		.h2f_rst_n                 (arria10_hps_0_h2f_reset_reset),                         //           h2f_reset.reset_n
		.f2h_cold_rst_req_n        (f2h_cold_reset_req_reset_n),                            //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n         (f2h_debug_reset_req_reset_n),                           // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n        (f2h_warm_reset_req_reset_n),                            //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents          (f2h_stm_hw_events_stm_hwevents),                        //   f2h_stm_hw_events.stm_hwevents
		.emif_emif_to_hps          (emif_a10_hps_0_hps_emif_conduit_end_emif_to_hps),       //                emif.emif_to_hps
		.emif_hps_to_emif          (arria10_hps_0_emif_hps_to_emif),                        //                    .hps_to_emif
		.emif_emif_to_gp           (emif_a10_hps_0_hps_emif_conduit_end_emif_to_gp),        //                    .emif_to_gp
		.emif_gp_to_emif           (arria10_hps_0_emif_gp_to_emif),                         //                    .gp_to_emif
		.f2h_axi_clk               (clk_100_clk),                                           //       f2h_axi_clock.clk
		.f2h_axi_rst               (~hps_fpga_reset_reset),                                 //       f2h_axi_reset.reset_n
		.f2h_AWID                  (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awid),    //       f2h_axi_slave.awid
		.f2h_AWADDR                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.f2h_AWLEN                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.f2h_AWSIZE                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.f2h_AWBURST               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.f2h_AWLOCK                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.f2h_AWCACHE               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.f2h_AWPROT                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.f2h_AWVALID               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.f2h_AWREADY               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awready), //                    .awready
		.f2h_AWUSER                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.f2h_WID                   (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wid),     //                    .wid
		.f2h_WDATA                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.f2h_WSTRB                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.f2h_WLAST                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.f2h_WVALID                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.f2h_WREADY                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wready),  //                    .wready
		.f2h_BID                   (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bid),     //                    .bid
		.f2h_BRESP                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.f2h_BVALID                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.f2h_BREADY                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bready),  //                    .bready
		.f2h_ARID                  (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arid),    //                    .arid
		.f2h_ARADDR                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.f2h_ARLEN                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.f2h_ARSIZE                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.f2h_ARBURST               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.f2h_ARLOCK                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.f2h_ARCACHE               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.f2h_ARPROT                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.f2h_ARVALID               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.f2h_ARREADY               (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arready), //                    .arready
		.f2h_ARUSER                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.f2h_RID                   (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rid),     //                    .rid
		.f2h_RDATA                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.f2h_RRESP                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.f2h_RLAST                 (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.f2h_RVALID                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.f2h_RREADY                (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rready),  //                    .rready
		.h2f_lw_axi_clk            (clk_100_clk),                                           //    h2f_lw_axi_clock.clk
		.h2f_lw_axi_rst            (~hps_fpga_reset_reset),                                 //    h2f_lw_axi_reset.reset_n
		.h2f_lw_AWID               (arria10_hps_0_h2f_lw_axi_master_awid),                  //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR             (arria10_hps_0_h2f_lw_axi_master_awaddr),                //                    .awaddr
		.h2f_lw_AWLEN              (arria10_hps_0_h2f_lw_axi_master_awlen),                 //                    .awlen
		.h2f_lw_AWSIZE             (arria10_hps_0_h2f_lw_axi_master_awsize),                //                    .awsize
		.h2f_lw_AWBURST            (arria10_hps_0_h2f_lw_axi_master_awburst),               //                    .awburst
		.h2f_lw_AWLOCK             (arria10_hps_0_h2f_lw_axi_master_awlock),                //                    .awlock
		.h2f_lw_AWCACHE            (arria10_hps_0_h2f_lw_axi_master_awcache),               //                    .awcache
		.h2f_lw_AWPROT             (arria10_hps_0_h2f_lw_axi_master_awprot),                //                    .awprot
		.h2f_lw_AWVALID            (arria10_hps_0_h2f_lw_axi_master_awvalid),               //                    .awvalid
		.h2f_lw_AWREADY            (arria10_hps_0_h2f_lw_axi_master_awready),               //                    .awready
		.h2f_lw_AWUSER             (arria10_hps_0_h2f_lw_axi_master_awuser),                //                    .awuser
		.h2f_lw_WID                (arria10_hps_0_h2f_lw_axi_master_wid),                   //                    .wid
		.h2f_lw_WDATA              (arria10_hps_0_h2f_lw_axi_master_wdata),                 //                    .wdata
		.h2f_lw_WSTRB              (arria10_hps_0_h2f_lw_axi_master_wstrb),                 //                    .wstrb
		.h2f_lw_WLAST              (arria10_hps_0_h2f_lw_axi_master_wlast),                 //                    .wlast
		.h2f_lw_WVALID             (arria10_hps_0_h2f_lw_axi_master_wvalid),                //                    .wvalid
		.h2f_lw_WREADY             (arria10_hps_0_h2f_lw_axi_master_wready),                //                    .wready
		.h2f_lw_BID                (arria10_hps_0_h2f_lw_axi_master_bid),                   //                    .bid
		.h2f_lw_BRESP              (arria10_hps_0_h2f_lw_axi_master_bresp),                 //                    .bresp
		.h2f_lw_BVALID             (arria10_hps_0_h2f_lw_axi_master_bvalid),                //                    .bvalid
		.h2f_lw_BREADY             (arria10_hps_0_h2f_lw_axi_master_bready),                //                    .bready
		.h2f_lw_ARID               (arria10_hps_0_h2f_lw_axi_master_arid),                  //                    .arid
		.h2f_lw_ARADDR             (arria10_hps_0_h2f_lw_axi_master_araddr),                //                    .araddr
		.h2f_lw_ARLEN              (arria10_hps_0_h2f_lw_axi_master_arlen),                 //                    .arlen
		.h2f_lw_ARSIZE             (arria10_hps_0_h2f_lw_axi_master_arsize),                //                    .arsize
		.h2f_lw_ARBURST            (arria10_hps_0_h2f_lw_axi_master_arburst),               //                    .arburst
		.h2f_lw_ARLOCK             (arria10_hps_0_h2f_lw_axi_master_arlock),                //                    .arlock
		.h2f_lw_ARCACHE            (arria10_hps_0_h2f_lw_axi_master_arcache),               //                    .arcache
		.h2f_lw_ARPROT             (arria10_hps_0_h2f_lw_axi_master_arprot),                //                    .arprot
		.h2f_lw_ARVALID            (arria10_hps_0_h2f_lw_axi_master_arvalid),               //                    .arvalid
		.h2f_lw_ARREADY            (arria10_hps_0_h2f_lw_axi_master_arready),               //                    .arready
		.h2f_lw_ARUSER             (arria10_hps_0_h2f_lw_axi_master_aruser),                //                    .aruser
		.h2f_lw_RID                (arria10_hps_0_h2f_lw_axi_master_rid),                   //                    .rid
		.h2f_lw_RDATA              (arria10_hps_0_h2f_lw_axi_master_rdata),                 //                    .rdata
		.h2f_lw_RRESP              (arria10_hps_0_h2f_lw_axi_master_rresp),                 //                    .rresp
		.h2f_lw_RLAST              (arria10_hps_0_h2f_lw_axi_master_rlast),                 //                    .rlast
		.h2f_lw_RVALID             (arria10_hps_0_h2f_lw_axi_master_rvalid),                //                    .rvalid
		.h2f_lw_RREADY             (arria10_hps_0_h2f_lw_axi_master_rready),                //                    .rready
		.h2f_axi_clk               (clk_100_clk),                                           //       h2f_axi_clock.clk
		.h2f_axi_rst               (~hps_fpga_reset_reset),                                 //       h2f_axi_reset.reset_n
		.h2f_AWID                  (arria10_hps_0_h2f_axi_master_awid),                     //      h2f_axi_master.awid
		.h2f_AWADDR                (arria10_hps_0_h2f_axi_master_awaddr),                   //                    .awaddr
		.h2f_AWLEN                 (arria10_hps_0_h2f_axi_master_awlen),                    //                    .awlen
		.h2f_AWSIZE                (arria10_hps_0_h2f_axi_master_awsize),                   //                    .awsize
		.h2f_AWBURST               (arria10_hps_0_h2f_axi_master_awburst),                  //                    .awburst
		.h2f_AWLOCK                (arria10_hps_0_h2f_axi_master_awlock),                   //                    .awlock
		.h2f_AWCACHE               (arria10_hps_0_h2f_axi_master_awcache),                  //                    .awcache
		.h2f_AWPROT                (arria10_hps_0_h2f_axi_master_awprot),                   //                    .awprot
		.h2f_AWVALID               (arria10_hps_0_h2f_axi_master_awvalid),                  //                    .awvalid
		.h2f_AWREADY               (arria10_hps_0_h2f_axi_master_awready),                  //                    .awready
		.h2f_AWUSER                (arria10_hps_0_h2f_axi_master_awuser),                   //                    .awuser
		.h2f_WID                   (arria10_hps_0_h2f_axi_master_wid),                      //                    .wid
		.h2f_WDATA                 (arria10_hps_0_h2f_axi_master_wdata),                    //                    .wdata
		.h2f_WSTRB                 (arria10_hps_0_h2f_axi_master_wstrb),                    //                    .wstrb
		.h2f_WLAST                 (arria10_hps_0_h2f_axi_master_wlast),                    //                    .wlast
		.h2f_WVALID                (arria10_hps_0_h2f_axi_master_wvalid),                   //                    .wvalid
		.h2f_WREADY                (arria10_hps_0_h2f_axi_master_wready),                   //                    .wready
		.h2f_BID                   (arria10_hps_0_h2f_axi_master_bid),                      //                    .bid
		.h2f_BRESP                 (arria10_hps_0_h2f_axi_master_bresp),                    //                    .bresp
		.h2f_BVALID                (arria10_hps_0_h2f_axi_master_bvalid),                   //                    .bvalid
		.h2f_BREADY                (arria10_hps_0_h2f_axi_master_bready),                   //                    .bready
		.h2f_ARID                  (arria10_hps_0_h2f_axi_master_arid),                     //                    .arid
		.h2f_ARADDR                (arria10_hps_0_h2f_axi_master_araddr),                   //                    .araddr
		.h2f_ARLEN                 (arria10_hps_0_h2f_axi_master_arlen),                    //                    .arlen
		.h2f_ARSIZE                (arria10_hps_0_h2f_axi_master_arsize),                   //                    .arsize
		.h2f_ARBURST               (arria10_hps_0_h2f_axi_master_arburst),                  //                    .arburst
		.h2f_ARLOCK                (arria10_hps_0_h2f_axi_master_arlock),                   //                    .arlock
		.h2f_ARCACHE               (arria10_hps_0_h2f_axi_master_arcache),                  //                    .arcache
		.h2f_ARPROT                (arria10_hps_0_h2f_axi_master_arprot),                   //                    .arprot
		.h2f_ARVALID               (arria10_hps_0_h2f_axi_master_arvalid),                  //                    .arvalid
		.h2f_ARREADY               (arria10_hps_0_h2f_axi_master_arready),                  //                    .arready
		.h2f_ARUSER                (arria10_hps_0_h2f_axi_master_aruser),                   //                    .aruser
		.h2f_RID                   (arria10_hps_0_h2f_axi_master_rid),                      //                    .rid
		.h2f_RDATA                 (arria10_hps_0_h2f_axi_master_rdata),                    //                    .rdata
		.h2f_RRESP                 (arria10_hps_0_h2f_axi_master_rresp),                    //                    .rresp
		.h2f_RLAST                 (arria10_hps_0_h2f_axi_master_rlast),                    //                    .rlast
		.h2f_RVALID                (arria10_hps_0_h2f_axi_master_rvalid),                   //                    .rvalid
		.h2f_RREADY                (arria10_hps_0_h2f_axi_master_rready),                   //                    .rready
		.f2sdram0_clk              (clk_100_clk),                                           //      f2sdram0_clock.clk
		.f2s_sdram0_rst            (~hps_fpga_reset_reset),                                 //      f2sdram0_reset.reset_n
		.f2sdram0_ARADDR           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_araddr),  //       f2sdram0_data.araddr
		.f2sdram0_ARBURST          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arburst), //                    .arburst
		.f2sdram0_ARCACHE          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arcache), //                    .arcache
		.f2sdram0_ARID             (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arid),    //                    .arid
		.f2sdram0_ARLEN            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlen),   //                    .arlen
		.f2sdram0_ARLOCK           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlock),  //                    .arlock
		.f2sdram0_ARPROT           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arprot),  //                    .arprot
		.f2sdram0_ARREADY          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arready), //                    .arready
		.f2sdram0_ARSIZE           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arsize),  //                    .arsize
		.f2sdram0_ARUSER           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_aruser),  //                    .aruser
		.f2sdram0_ARVALID          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arvalid), //                    .arvalid
		.f2sdram0_AWADDR           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awaddr),  //                    .awaddr
		.f2sdram0_AWBURST          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awburst), //                    .awburst
		.f2sdram0_AWCACHE          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awcache), //                    .awcache
		.f2sdram0_AWID             (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awid),    //                    .awid
		.f2sdram0_AWLEN            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlen),   //                    .awlen
		.f2sdram0_AWLOCK           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlock),  //                    .awlock
		.f2sdram0_AWPROT           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awprot),  //                    .awprot
		.f2sdram0_AWREADY          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awready), //                    .awready
		.f2sdram0_AWSIZE           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awsize),  //                    .awsize
		.f2sdram0_AWUSER           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awuser),  //                    .awuser
		.f2sdram0_AWVALID          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awvalid), //                    .awvalid
		.f2sdram0_WDATA            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wdata),   //                    .wdata
		.f2sdram0_WID              (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wid),     //                    .wid
		.f2sdram0_WLAST            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wlast),   //                    .wlast
		.f2sdram0_WREADY           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wready),  //                    .wready
		.f2sdram0_WSTRB            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wstrb),   //                    .wstrb
		.f2sdram0_WVALID           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wvalid),  //                    .wvalid
		.f2sdram0_BID              (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bid),     //                    .bid
		.f2sdram0_BREADY           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bready),  //                    .bready
		.f2sdram0_BRESP            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bresp),   //                    .bresp
		.f2sdram0_BVALID           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bvalid),  //                    .bvalid
		.f2sdram0_RDATA            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rdata),   //                    .rdata
		.f2sdram0_RID              (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rid),     //                    .rid
		.f2sdram0_RLAST            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rlast),   //                    .rlast
		.f2sdram0_RREADY           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rready),  //                    .rready
		.f2sdram0_RRESP            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rresp),   //                    .rresp
		.f2sdram0_RVALID           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rvalid),  //                    .rvalid
		.f2sdram2_clk              (clk_100_clk),                                           //      f2sdram2_clock.clk
		.f2s_sdram2_rst            (~hps_fpga_reset_reset),                                 //      f2sdram2_reset.reset_n
		.f2sdram2_ARADDR           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_araddr),  //       f2sdram2_data.araddr
		.f2sdram2_ARBURST          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arburst), //                    .arburst
		.f2sdram2_ARCACHE          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arcache), //                    .arcache
		.f2sdram2_ARID             (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arid),    //                    .arid
		.f2sdram2_ARLEN            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlen),   //                    .arlen
		.f2sdram2_ARLOCK           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlock),  //                    .arlock
		.f2sdram2_ARPROT           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arprot),  //                    .arprot
		.f2sdram2_ARREADY          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arready), //                    .arready
		.f2sdram2_ARSIZE           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arsize),  //                    .arsize
		.f2sdram2_ARUSER           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_aruser),  //                    .aruser
		.f2sdram2_ARVALID          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arvalid), //                    .arvalid
		.f2sdram2_AWADDR           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awaddr),  //                    .awaddr
		.f2sdram2_AWBURST          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awburst), //                    .awburst
		.f2sdram2_AWCACHE          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awcache), //                    .awcache
		.f2sdram2_AWID             (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awid),    //                    .awid
		.f2sdram2_AWLEN            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlen),   //                    .awlen
		.f2sdram2_AWLOCK           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlock),  //                    .awlock
		.f2sdram2_AWPROT           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awprot),  //                    .awprot
		.f2sdram2_AWREADY          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awready), //                    .awready
		.f2sdram2_AWSIZE           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awsize),  //                    .awsize
		.f2sdram2_AWUSER           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awuser),  //                    .awuser
		.f2sdram2_AWVALID          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awvalid), //                    .awvalid
		.f2sdram2_WDATA            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wdata),   //                    .wdata
		.f2sdram2_WID              (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wid),     //                    .wid
		.f2sdram2_WLAST            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wlast),   //                    .wlast
		.f2sdram2_WREADY           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wready),  //                    .wready
		.f2sdram2_WSTRB            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wstrb),   //                    .wstrb
		.f2sdram2_WVALID           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wvalid),  //                    .wvalid
		.f2sdram2_BID              (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bid),     //                    .bid
		.f2sdram2_BREADY           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bready),  //                    .bready
		.f2sdram2_BRESP            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bresp),   //                    .bresp
		.f2sdram2_BVALID           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bvalid),  //                    .bvalid
		.f2sdram2_RDATA            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rdata),   //                    .rdata
		.f2sdram2_RID              (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rid),     //                    .rid
		.f2sdram2_RLAST            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rlast),   //                    .rlast
		.f2sdram2_RREADY           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rready),  //                    .rready
		.f2sdram2_RRESP            (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rresp),   //                    .rresp
		.f2sdram2_RVALID           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rvalid),  //                    .rvalid
		.f2h_irq_p0                (arria10_hps_0_f2h_irq0_irq),                            //            f2h_irq0.irq
		.f2h_irq_p1                (arria10_hps_0_f2h_irq1_irq),                            //            f2h_irq1.irq
		.hps_io_phery_emac0_TX_CLK (hps_io_hps_io_phery_emac0_TX_CLK),                      //              hps_io.hps_io_phery_emac0_TX_CLK
		.hps_io_phery_emac0_TXD0   (hps_io_hps_io_phery_emac0_TXD0),                        //                    .hps_io_phery_emac0_TXD0
		.hps_io_phery_emac0_TXD1   (hps_io_hps_io_phery_emac0_TXD1),                        //                    .hps_io_phery_emac0_TXD1
		.hps_io_phery_emac0_TXD2   (hps_io_hps_io_phery_emac0_TXD2),                        //                    .hps_io_phery_emac0_TXD2
		.hps_io_phery_emac0_TXD3   (hps_io_hps_io_phery_emac0_TXD3),                        //                    .hps_io_phery_emac0_TXD3
		.hps_io_phery_emac0_RX_CTL (hps_io_hps_io_phery_emac0_RX_CTL),                      //                    .hps_io_phery_emac0_RX_CTL
		.hps_io_phery_emac0_TX_CTL (hps_io_hps_io_phery_emac0_TX_CTL),                      //                    .hps_io_phery_emac0_TX_CTL
		.hps_io_phery_emac0_RX_CLK (hps_io_hps_io_phery_emac0_RX_CLK),                      //                    .hps_io_phery_emac0_RX_CLK
		.hps_io_phery_emac0_RXD0   (hps_io_hps_io_phery_emac0_RXD0),                        //                    .hps_io_phery_emac0_RXD0
		.hps_io_phery_emac0_RXD1   (hps_io_hps_io_phery_emac0_RXD1),                        //                    .hps_io_phery_emac0_RXD1
		.hps_io_phery_emac0_RXD2   (hps_io_hps_io_phery_emac0_RXD2),                        //                    .hps_io_phery_emac0_RXD2
		.hps_io_phery_emac0_RXD3   (hps_io_hps_io_phery_emac0_RXD3),                        //                    .hps_io_phery_emac0_RXD3
		.hps_io_phery_emac0_MDIO   (hps_io_hps_io_phery_emac0_MDIO),                        //                    .hps_io_phery_emac0_MDIO
		.hps_io_phery_emac0_MDC    (hps_io_hps_io_phery_emac0_MDC),                         //                    .hps_io_phery_emac0_MDC
		.hps_io_phery_sdmmc_CMD    (hps_io_hps_io_phery_sdmmc_CMD),                         //                    .hps_io_phery_sdmmc_CMD
		.hps_io_phery_sdmmc_D0     (hps_io_hps_io_phery_sdmmc_D0),                          //                    .hps_io_phery_sdmmc_D0
		.hps_io_phery_sdmmc_D1     (hps_io_hps_io_phery_sdmmc_D1),                          //                    .hps_io_phery_sdmmc_D1
		.hps_io_phery_sdmmc_D2     (hps_io_hps_io_phery_sdmmc_D2),                          //                    .hps_io_phery_sdmmc_D2
		.hps_io_phery_sdmmc_D3     (hps_io_hps_io_phery_sdmmc_D3),                          //                    .hps_io_phery_sdmmc_D3
		.hps_io_phery_sdmmc_D4     (hps_io_hps_io_phery_sdmmc_D4),                          //                    .hps_io_phery_sdmmc_D4
		.hps_io_phery_sdmmc_D5     (hps_io_hps_io_phery_sdmmc_D5),                          //                    .hps_io_phery_sdmmc_D5
		.hps_io_phery_sdmmc_D6     (hps_io_hps_io_phery_sdmmc_D6),                          //                    .hps_io_phery_sdmmc_D6
		.hps_io_phery_sdmmc_D7     (hps_io_hps_io_phery_sdmmc_D7),                          //                    .hps_io_phery_sdmmc_D7
		.hps_io_phery_sdmmc_CCLK   (hps_io_hps_io_phery_sdmmc_CCLK),                        //                    .hps_io_phery_sdmmc_CCLK
		.hps_io_phery_usb0_DATA0   (hps_io_hps_io_phery_usb0_DATA0),                        //                    .hps_io_phery_usb0_DATA0
		.hps_io_phery_usb0_DATA1   (hps_io_hps_io_phery_usb0_DATA1),                        //                    .hps_io_phery_usb0_DATA1
		.hps_io_phery_usb0_DATA2   (hps_io_hps_io_phery_usb0_DATA2),                        //                    .hps_io_phery_usb0_DATA2
		.hps_io_phery_usb0_DATA3   (hps_io_hps_io_phery_usb0_DATA3),                        //                    .hps_io_phery_usb0_DATA3
		.hps_io_phery_usb0_DATA4   (hps_io_hps_io_phery_usb0_DATA4),                        //                    .hps_io_phery_usb0_DATA4
		.hps_io_phery_usb0_DATA5   (hps_io_hps_io_phery_usb0_DATA5),                        //                    .hps_io_phery_usb0_DATA5
		.hps_io_phery_usb0_DATA6   (hps_io_hps_io_phery_usb0_DATA6),                        //                    .hps_io_phery_usb0_DATA6
		.hps_io_phery_usb0_DATA7   (hps_io_hps_io_phery_usb0_DATA7),                        //                    .hps_io_phery_usb0_DATA7
		.hps_io_phery_usb0_CLK     (hps_io_hps_io_phery_usb0_CLK),                          //                    .hps_io_phery_usb0_CLK
		.hps_io_phery_usb0_STP     (hps_io_hps_io_phery_usb0_STP),                          //                    .hps_io_phery_usb0_STP
		.hps_io_phery_usb0_DIR     (hps_io_hps_io_phery_usb0_DIR),                          //                    .hps_io_phery_usb0_DIR
		.hps_io_phery_usb0_NXT     (hps_io_hps_io_phery_usb0_NXT),                          //                    .hps_io_phery_usb0_NXT
		.hps_io_phery_spim1_CLK    (hps_io_hps_io_phery_spim1_CLK),                         //                    .hps_io_phery_spim1_CLK
		.hps_io_phery_spim1_MOSI   (hps_io_hps_io_phery_spim1_MOSI),                        //                    .hps_io_phery_spim1_MOSI
		.hps_io_phery_spim1_MISO   (hps_io_hps_io_phery_spim1_MISO),                        //                    .hps_io_phery_spim1_MISO
		.hps_io_phery_spim1_SS0_N  (hps_io_hps_io_phery_spim1_SS0_N),                       //                    .hps_io_phery_spim1_SS0_N
		.hps_io_phery_spim1_SS1_N  (hps_io_hps_io_phery_spim1_SS1_N),                       //                    .hps_io_phery_spim1_SS1_N
		.hps_io_phery_trace_CLK    (hps_io_hps_io_phery_trace_CLK),                         //                    .hps_io_phery_trace_CLK
		.hps_io_phery_trace_D0     (hps_io_hps_io_phery_trace_D0),                          //                    .hps_io_phery_trace_D0
		.hps_io_phery_trace_D1     (hps_io_hps_io_phery_trace_D1),                          //                    .hps_io_phery_trace_D1
		.hps_io_phery_trace_D2     (hps_io_hps_io_phery_trace_D2),                          //                    .hps_io_phery_trace_D2
		.hps_io_phery_trace_D3     (hps_io_hps_io_phery_trace_D3),                          //                    .hps_io_phery_trace_D3
		.hps_io_phery_uart1_RX     (hps_io_hps_io_phery_uart1_RX),                          //                    .hps_io_phery_uart1_RX
		.hps_io_phery_uart1_TX     (hps_io_hps_io_phery_uart1_TX),                          //                    .hps_io_phery_uart1_TX
		.hps_io_phery_i2c1_SDA     (hps_io_hps_io_phery_i2c1_SDA),                          //                    .hps_io_phery_i2c1_SDA
		.hps_io_phery_i2c1_SCL     (hps_io_hps_io_phery_i2c1_SCL),                          //                    .hps_io_phery_i2c1_SCL
		.hps_io_gpio_gpio1_io5     (hps_io_hps_io_gpio_gpio1_io5),                          //                    .hps_io_gpio_gpio1_io5
		.hps_io_gpio_gpio1_io14    (hps_io_hps_io_gpio_gpio1_io14),                         //                    .hps_io_gpio_gpio1_io14
		.hps_io_gpio_gpio1_io16    (hps_io_hps_io_gpio_gpio1_io16),                         //                    .hps_io_gpio_gpio1_io16
		.hps_io_gpio_gpio1_io17    (hps_io_hps_io_gpio_gpio1_io17)                          //                    .hps_io_gpio_gpio1_io17
	);

	ghrd_10as066n2_altera_avalon_pio_161_imbvr3i button_pio (
		.clk        (clk_100_clk),                                //                 clk.clk
		.reset_n    (~hps_fpga_reset_reset),                      //               reset.reset_n
		.address    (mm_interconnect_2_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_button_pio_s1_readdata),   //                    .readdata
		.in_port    (pio_button_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                    //                 irq.irq
	);

	ghrd_10as066n2_altera_avalon_pio_161_wd25eay dipsw_pio (
		.clk        (clk_100_clk),                               //                 clk.clk
		.reset_n    (~hps_fpga_reset_reset),                     //               reset.reset_n
		.address    (mm_interconnect_2_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_dipsw_pio_s1_readdata),   //                    .readdata
		.in_port    (pio_dipsw_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	ghrd_10as066n2_altera_emif_a10_hps_161_6mh7udq emif_a10_hps_0 (
		.global_reset_n (reset_reset_n),                                   // global_reset_reset_sink.reset_n
		.pll_ref_clk    (emif_a10_hps_0_pll_ref_clk_clock_sink_clk),       //  pll_ref_clk_clock_sink.clk
		.oct_rzqin      (emif_a10_hps_0_oct_conduit_end_oct_rzqin),        //         oct_conduit_end.oct_rzqin
		.mem_ck         (emif_a10_hps_0_mem_conduit_end_mem_ck),           //         mem_conduit_end.mem_ck
		.mem_ck_n       (emif_a10_hps_0_mem_conduit_end_mem_ck_n),         //                        .mem_ck_n
		.mem_a          (emif_a10_hps_0_mem_conduit_end_mem_a),            //                        .mem_a
		.mem_act_n      (emif_a10_hps_0_mem_conduit_end_mem_act_n),        //                        .mem_act_n
		.mem_ba         (emif_a10_hps_0_mem_conduit_end_mem_ba),           //                        .mem_ba
		.mem_bg         (emif_a10_hps_0_mem_conduit_end_mem_bg),           //                        .mem_bg
		.mem_cke        (emif_a10_hps_0_mem_conduit_end_mem_cke),          //                        .mem_cke
		.mem_cs_n       (emif_a10_hps_0_mem_conduit_end_mem_cs_n),         //                        .mem_cs_n
		.mem_odt        (emif_a10_hps_0_mem_conduit_end_mem_odt),          //                        .mem_odt
		.mem_reset_n    (emif_a10_hps_0_mem_conduit_end_mem_reset_n),      //                        .mem_reset_n
		.mem_par        (emif_a10_hps_0_mem_conduit_end_mem_par),          //                        .mem_par
		.mem_alert_n    (emif_a10_hps_0_mem_conduit_end_mem_alert_n),      //                        .mem_alert_n
		.mem_dqs        (emif_a10_hps_0_mem_conduit_end_mem_dqs),          //                        .mem_dqs
		.mem_dqs_n      (emif_a10_hps_0_mem_conduit_end_mem_dqs_n),        //                        .mem_dqs_n
		.mem_dq         (emif_a10_hps_0_mem_conduit_end_mem_dq),           //                        .mem_dq
		.mem_dbi_n      (emif_a10_hps_0_mem_conduit_end_mem_dbi_n),        //                        .mem_dbi_n
		.hps_to_emif    (arria10_hps_0_emif_hps_to_emif),                  //    hps_emif_conduit_end.hps_to_emif
		.emif_to_hps    (emif_a10_hps_0_hps_emif_conduit_end_emif_to_hps), //                        .emif_to_hps
		.hps_to_emif_gp (arria10_hps_0_emif_gp_to_emif),                   //                        .gp_to_emif
		.emif_to_hps_gp (emif_a10_hps_0_hps_emif_conduit_end_emif_to_gp)   //                        .emif_to_gp
	);

	ghrd_10as066n2_altera_jtag_avalon_master_161_7opu3yi #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) f2sdram_only_master (
		.clk_clk              (clk_100_clk),                              //          clk.clk
		.clk_reset_reset      (rst_controller_001_reset_out_reset),       //    clk_reset.reset
		.master_address       (f2sdram_only_master_master_address),       //       master.address
		.master_readdata      (f2sdram_only_master_master_readdata),      //             .readdata
		.master_read          (f2sdram_only_master_master_read),          //             .read
		.master_write         (f2sdram_only_master_master_write),         //             .write
		.master_writedata     (f2sdram_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (f2sdram_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (f2sdram_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (f2sdram_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	ghrd_10as066n2_altera_jtag_avalon_master_161_7opu3yi #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) f2sdram_only_master1 (
		.clk_clk              (clk_100_clk),                               //          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset),        //    clk_reset.reset
		.master_address       (f2sdram_only_master1_master_address),       //       master.address
		.master_readdata      (f2sdram_only_master1_master_readdata),      //             .readdata
		.master_read          (f2sdram_only_master1_master_read),          //             .read
		.master_write         (f2sdram_only_master1_master_write),         //             .write
		.master_writedata     (f2sdram_only_master1_master_writedata),     //             .writedata
		.master_waitrequest   (f2sdram_only_master1_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (f2sdram_only_master1_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (f2sdram_only_master1_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                           // master_reset.reset
	);

	ghrd_10as066n2_altera_jtag_avalon_master_161_7opu3yi #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (clk_100_clk),                           //          clk.clk
		.clk_reset_reset      (rst_controller_003_reset_out_reset),    //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	ghrd_10as066n2_altera_jtag_avalon_master_161_7opu3yi #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_only_master (
		.clk_clk              (clk_100_clk),                          //          clk.clk
		.clk_reset_reset      (rst_controller_004_reset_out_reset),   //    clk_reset.reset
		.master_address       (hps_only_master_master_address),       //       master.address
		.master_readdata      (hps_only_master_master_readdata),      //             .readdata
		.master_read          (hps_only_master_master_read),          //             .read
		.master_write         (hps_only_master_master_write),         //             .write
		.master_writedata     (hps_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                      // master_reset.reset
	);

	altsource_probe #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("RST"),
		.probe_width             (0),
		.source_width            (3),
		.source_initial_value    ("0"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (issp_hps_resets_source), //    sources.source
		.source_clk (clk_100_clk),            // source_clk.clk
		.source_ena (1'b1)                    // (terminated)
	);

	ghrd_10as066n2_altera_avalon_pio_161_p5oy5va led_pio (
		.clk        (clk_100_clk),                             //                 clk.clk
		.reset_n    (~hps_fpga_reset_reset),                   //               reset.reset_n
		.address    (mm_interconnect_2_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_led_pio_s1_readdata),   //                    .readdata
		.in_port    (pio_led_external_connection_in_port),     // external_connection.export
		.out_port   (pio_led_external_connection_out_port)     //                    .export
	);

	ghrd_10as066n2_altera_avalon_onchip_memory2_161_lxrufkq onchip_memory2_0 (
		.clk        (clk_100_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.reset      (hps_fpga_reset_reset),                             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (9),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pb_lwh2f (
		.clk              (clk_100_clk),                                 //   clk.clk
		.reset            (hps_fpga_reset_reset),                        // reset.reset
		.s0_waitrequest   (mm_interconnect_1_pb_lwh2f_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_pb_lwh2f_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_pb_lwh2f_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_pb_lwh2f_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_pb_lwh2f_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_pb_lwh2f_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_pb_lwh2f_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_pb_lwh2f_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_pb_lwh2f_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_pb_lwh2f_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pb_lwh2f_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pb_lwh2f_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pb_lwh2f_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pb_lwh2f_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pb_lwh2f_m0_writedata),                       //      .writedata
		.m0_address       (pb_lwh2f_m0_address),                         //      .address
		.m0_write         (pb_lwh2f_m0_write),                           //      .write
		.m0_read          (pb_lwh2f_m0_read),                            //      .read
		.m0_byteenable    (pb_lwh2f_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pb_lwh2f_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                            // (terminated)
		.m0_response      (2'b00)                                        // (terminated)
	);

	protobuf_serializer protobuf_serializer_0 (
		.clock_clk      (clk_100_clk),                                        // clock.clk
		.reset_reset_n  (~hps_fpga_reset_reset),                              // reset.reset_n
		.axs_s0_wstrb   (mm_interconnect_0_protobuf_serializer_0_s0_wstrb),   //    s0.wstrb
		.axs_s0_wready  (mm_interconnect_0_protobuf_serializer_0_s0_wready),  //      .wready
		.axs_s0_wdata   (mm_interconnect_0_protobuf_serializer_0_s0_wdata),   //      .wdata
		.axs_s0_rvalid  (mm_interconnect_0_protobuf_serializer_0_s0_rvalid),  //      .rvalid
		.axs_s0_rready  (mm_interconnect_0_protobuf_serializer_0_s0_rready),  //      .rready
		.axs_s0_rlast   (mm_interconnect_0_protobuf_serializer_0_s0_rlast),   //      .rlast
		.axs_s0_rid     (mm_interconnect_0_protobuf_serializer_0_s0_rid),     //      .rid
		.axs_s0_rdata   (mm_interconnect_0_protobuf_serializer_0_s0_rdata),   //      .rdata
		.axs_s0_bvalid  (mm_interconnect_0_protobuf_serializer_0_s0_bvalid),  //      .bvalid
		.axs_s0_bready  (mm_interconnect_0_protobuf_serializer_0_s0_bready),  //      .bready
		.axs_s0_bid     (mm_interconnect_0_protobuf_serializer_0_s0_bid),     //      .bid
		.axs_s0_awsize  (mm_interconnect_0_protobuf_serializer_0_s0_awsize),  //      .awsize
		.axs_s0_awready (mm_interconnect_0_protobuf_serializer_0_s0_awready), //      .awready
		.axs_s0_awlen   (mm_interconnect_0_protobuf_serializer_0_s0_awlen),   //      .awlen
		.axs_s0_awid    (mm_interconnect_0_protobuf_serializer_0_s0_awid),    //      .awid
		.axs_s0_awburst (mm_interconnect_0_protobuf_serializer_0_s0_awburst), //      .awburst
		.axs_s0_awaddr  (mm_interconnect_0_protobuf_serializer_0_s0_awaddr),  //      .awaddr
		.axs_s0_arvalid (mm_interconnect_0_protobuf_serializer_0_s0_arvalid), //      .arvalid
		.axs_s0_arsize  (mm_interconnect_0_protobuf_serializer_0_s0_arsize),  //      .arsize
		.axs_s0_arready (mm_interconnect_0_protobuf_serializer_0_s0_arready), //      .arready
		.axs_s0_arlen   (mm_interconnect_0_protobuf_serializer_0_s0_arlen),   //      .arlen
		.axs_s0_arid    (mm_interconnect_0_protobuf_serializer_0_s0_arid),    //      .arid
		.axs_s0_arburst (mm_interconnect_0_protobuf_serializer_0_s0_arburst), //      .arburst
		.axs_s0_araddr  (mm_interconnect_0_protobuf_serializer_0_s0_araddr),  //      .araddr
		.axs_s0_wvalid  (mm_interconnect_0_protobuf_serializer_0_s0_wvalid),  //      .wvalid
		.axs_s0_awvalid (mm_interconnect_0_protobuf_serializer_0_s0_awvalid)  //      .awvalid
	);

	ghrd_10as066n2_altera_avalon_sysid_qsys_161_qri4vpa sysid_qsys_0 (
		.clock    (clk_100_clk),                                           //           clk.clk
		.reset_n  (~hps_fpga_reset_reset),                                 //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_0_control_slave_address)   //              .address
	);

	ghrd_10as066n2_altera_mm_interconnect_161_yundlma mm_interconnect_0 (
		.arria10_hps_0_h2f_axi_master_awid                       (arria10_hps_0_h2f_axi_master_awid),                  //                      arria10_hps_0_h2f_axi_master.awid
		.arria10_hps_0_h2f_axi_master_awaddr                     (arria10_hps_0_h2f_axi_master_awaddr),                //                                                  .awaddr
		.arria10_hps_0_h2f_axi_master_awlen                      (arria10_hps_0_h2f_axi_master_awlen),                 //                                                  .awlen
		.arria10_hps_0_h2f_axi_master_awsize                     (arria10_hps_0_h2f_axi_master_awsize),                //                                                  .awsize
		.arria10_hps_0_h2f_axi_master_awburst                    (arria10_hps_0_h2f_axi_master_awburst),               //                                                  .awburst
		.arria10_hps_0_h2f_axi_master_awlock                     (arria10_hps_0_h2f_axi_master_awlock),                //                                                  .awlock
		.arria10_hps_0_h2f_axi_master_awcache                    (arria10_hps_0_h2f_axi_master_awcache),               //                                                  .awcache
		.arria10_hps_0_h2f_axi_master_awprot                     (arria10_hps_0_h2f_axi_master_awprot),                //                                                  .awprot
		.arria10_hps_0_h2f_axi_master_awuser                     (arria10_hps_0_h2f_axi_master_awuser),                //                                                  .awuser
		.arria10_hps_0_h2f_axi_master_awvalid                    (arria10_hps_0_h2f_axi_master_awvalid),               //                                                  .awvalid
		.arria10_hps_0_h2f_axi_master_awready                    (arria10_hps_0_h2f_axi_master_awready),               //                                                  .awready
		.arria10_hps_0_h2f_axi_master_wid                        (arria10_hps_0_h2f_axi_master_wid),                   //                                                  .wid
		.arria10_hps_0_h2f_axi_master_wdata                      (arria10_hps_0_h2f_axi_master_wdata),                 //                                                  .wdata
		.arria10_hps_0_h2f_axi_master_wstrb                      (arria10_hps_0_h2f_axi_master_wstrb),                 //                                                  .wstrb
		.arria10_hps_0_h2f_axi_master_wlast                      (arria10_hps_0_h2f_axi_master_wlast),                 //                                                  .wlast
		.arria10_hps_0_h2f_axi_master_wvalid                     (arria10_hps_0_h2f_axi_master_wvalid),                //                                                  .wvalid
		.arria10_hps_0_h2f_axi_master_wready                     (arria10_hps_0_h2f_axi_master_wready),                //                                                  .wready
		.arria10_hps_0_h2f_axi_master_bid                        (arria10_hps_0_h2f_axi_master_bid),                   //                                                  .bid
		.arria10_hps_0_h2f_axi_master_bresp                      (arria10_hps_0_h2f_axi_master_bresp),                 //                                                  .bresp
		.arria10_hps_0_h2f_axi_master_bvalid                     (arria10_hps_0_h2f_axi_master_bvalid),                //                                                  .bvalid
		.arria10_hps_0_h2f_axi_master_bready                     (arria10_hps_0_h2f_axi_master_bready),                //                                                  .bready
		.arria10_hps_0_h2f_axi_master_arid                       (arria10_hps_0_h2f_axi_master_arid),                  //                                                  .arid
		.arria10_hps_0_h2f_axi_master_araddr                     (arria10_hps_0_h2f_axi_master_araddr),                //                                                  .araddr
		.arria10_hps_0_h2f_axi_master_arlen                      (arria10_hps_0_h2f_axi_master_arlen),                 //                                                  .arlen
		.arria10_hps_0_h2f_axi_master_arsize                     (arria10_hps_0_h2f_axi_master_arsize),                //                                                  .arsize
		.arria10_hps_0_h2f_axi_master_arburst                    (arria10_hps_0_h2f_axi_master_arburst),               //                                                  .arburst
		.arria10_hps_0_h2f_axi_master_arlock                     (arria10_hps_0_h2f_axi_master_arlock),                //                                                  .arlock
		.arria10_hps_0_h2f_axi_master_arcache                    (arria10_hps_0_h2f_axi_master_arcache),               //                                                  .arcache
		.arria10_hps_0_h2f_axi_master_arprot                     (arria10_hps_0_h2f_axi_master_arprot),                //                                                  .arprot
		.arria10_hps_0_h2f_axi_master_aruser                     (arria10_hps_0_h2f_axi_master_aruser),                //                                                  .aruser
		.arria10_hps_0_h2f_axi_master_arvalid                    (arria10_hps_0_h2f_axi_master_arvalid),               //                                                  .arvalid
		.arria10_hps_0_h2f_axi_master_arready                    (arria10_hps_0_h2f_axi_master_arready),               //                                                  .arready
		.arria10_hps_0_h2f_axi_master_rid                        (arria10_hps_0_h2f_axi_master_rid),                   //                                                  .rid
		.arria10_hps_0_h2f_axi_master_rdata                      (arria10_hps_0_h2f_axi_master_rdata),                 //                                                  .rdata
		.arria10_hps_0_h2f_axi_master_rresp                      (arria10_hps_0_h2f_axi_master_rresp),                 //                                                  .rresp
		.arria10_hps_0_h2f_axi_master_rlast                      (arria10_hps_0_h2f_axi_master_rlast),                 //                                                  .rlast
		.arria10_hps_0_h2f_axi_master_rvalid                     (arria10_hps_0_h2f_axi_master_rvalid),                //                                                  .rvalid
		.arria10_hps_0_h2f_axi_master_rready                     (arria10_hps_0_h2f_axi_master_rready),                //                                                  .rready
		.protobuf_serializer_0_s0_awid                           (mm_interconnect_0_protobuf_serializer_0_s0_awid),    //                          protobuf_serializer_0_s0.awid
		.protobuf_serializer_0_s0_awaddr                         (mm_interconnect_0_protobuf_serializer_0_s0_awaddr),  //                                                  .awaddr
		.protobuf_serializer_0_s0_awlen                          (mm_interconnect_0_protobuf_serializer_0_s0_awlen),   //                                                  .awlen
		.protobuf_serializer_0_s0_awsize                         (mm_interconnect_0_protobuf_serializer_0_s0_awsize),  //                                                  .awsize
		.protobuf_serializer_0_s0_awburst                        (mm_interconnect_0_protobuf_serializer_0_s0_awburst), //                                                  .awburst
		.protobuf_serializer_0_s0_awvalid                        (mm_interconnect_0_protobuf_serializer_0_s0_awvalid), //                                                  .awvalid
		.protobuf_serializer_0_s0_awready                        (mm_interconnect_0_protobuf_serializer_0_s0_awready), //                                                  .awready
		.protobuf_serializer_0_s0_wdata                          (mm_interconnect_0_protobuf_serializer_0_s0_wdata),   //                                                  .wdata
		.protobuf_serializer_0_s0_wstrb                          (mm_interconnect_0_protobuf_serializer_0_s0_wstrb),   //                                                  .wstrb
		.protobuf_serializer_0_s0_wvalid                         (mm_interconnect_0_protobuf_serializer_0_s0_wvalid),  //                                                  .wvalid
		.protobuf_serializer_0_s0_wready                         (mm_interconnect_0_protobuf_serializer_0_s0_wready),  //                                                  .wready
		.protobuf_serializer_0_s0_bid                            (mm_interconnect_0_protobuf_serializer_0_s0_bid),     //                                                  .bid
		.protobuf_serializer_0_s0_bvalid                         (mm_interconnect_0_protobuf_serializer_0_s0_bvalid),  //                                                  .bvalid
		.protobuf_serializer_0_s0_bready                         (mm_interconnect_0_protobuf_serializer_0_s0_bready),  //                                                  .bready
		.protobuf_serializer_0_s0_arid                           (mm_interconnect_0_protobuf_serializer_0_s0_arid),    //                                                  .arid
		.protobuf_serializer_0_s0_araddr                         (mm_interconnect_0_protobuf_serializer_0_s0_araddr),  //                                                  .araddr
		.protobuf_serializer_0_s0_arlen                          (mm_interconnect_0_protobuf_serializer_0_s0_arlen),   //                                                  .arlen
		.protobuf_serializer_0_s0_arsize                         (mm_interconnect_0_protobuf_serializer_0_s0_arsize),  //                                                  .arsize
		.protobuf_serializer_0_s0_arburst                        (mm_interconnect_0_protobuf_serializer_0_s0_arburst), //                                                  .arburst
		.protobuf_serializer_0_s0_arvalid                        (mm_interconnect_0_protobuf_serializer_0_s0_arvalid), //                                                  .arvalid
		.protobuf_serializer_0_s0_arready                        (mm_interconnect_0_protobuf_serializer_0_s0_arready), //                                                  .arready
		.protobuf_serializer_0_s0_rid                            (mm_interconnect_0_protobuf_serializer_0_s0_rid),     //                                                  .rid
		.protobuf_serializer_0_s0_rdata                          (mm_interconnect_0_protobuf_serializer_0_s0_rdata),   //                                                  .rdata
		.protobuf_serializer_0_s0_rlast                          (mm_interconnect_0_protobuf_serializer_0_s0_rlast),   //                                                  .rlast
		.protobuf_serializer_0_s0_rvalid                         (mm_interconnect_0_protobuf_serializer_0_s0_rvalid),  //                                                  .rvalid
		.protobuf_serializer_0_s0_rready                         (mm_interconnect_0_protobuf_serializer_0_s0_rready),  //                                                  .rready
		.clk_0_clk_clk                                           (clk_100_clk),                                        //                                         clk_0_clk.clk
		.arria10_hps_0_h2f_axi_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                               // arria10_hps_0_h2f_axi_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_s1_address                             (mm_interconnect_0_onchip_memory2_0_s1_address),      //                               onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                               (mm_interconnect_0_onchip_memory2_0_s1_write),        //                                                  .write
		.onchip_memory2_0_s1_readdata                            (mm_interconnect_0_onchip_memory2_0_s1_readdata),     //                                                  .readdata
		.onchip_memory2_0_s1_writedata                           (mm_interconnect_0_onchip_memory2_0_s1_writedata),    //                                                  .writedata
		.onchip_memory2_0_s1_chipselect                          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),   //                                                  .chipselect
		.onchip_memory2_0_s1_clken                               (mm_interconnect_0_onchip_memory2_0_s1_clken)         //                                                  .clken
	);

	ghrd_10as066n2_altera_mm_interconnect_161_k5z5r4y mm_interconnect_1 (
		.arria10_hps_0_h2f_lw_axi_master_awid                       (arria10_hps_0_h2f_lw_axi_master_awid),        //                      arria10_hps_0_h2f_lw_axi_master.awid
		.arria10_hps_0_h2f_lw_axi_master_awaddr                     (arria10_hps_0_h2f_lw_axi_master_awaddr),      //                                                     .awaddr
		.arria10_hps_0_h2f_lw_axi_master_awlen                      (arria10_hps_0_h2f_lw_axi_master_awlen),       //                                                     .awlen
		.arria10_hps_0_h2f_lw_axi_master_awsize                     (arria10_hps_0_h2f_lw_axi_master_awsize),      //                                                     .awsize
		.arria10_hps_0_h2f_lw_axi_master_awburst                    (arria10_hps_0_h2f_lw_axi_master_awburst),     //                                                     .awburst
		.arria10_hps_0_h2f_lw_axi_master_awlock                     (arria10_hps_0_h2f_lw_axi_master_awlock),      //                                                     .awlock
		.arria10_hps_0_h2f_lw_axi_master_awcache                    (arria10_hps_0_h2f_lw_axi_master_awcache),     //                                                     .awcache
		.arria10_hps_0_h2f_lw_axi_master_awprot                     (arria10_hps_0_h2f_lw_axi_master_awprot),      //                                                     .awprot
		.arria10_hps_0_h2f_lw_axi_master_awuser                     (arria10_hps_0_h2f_lw_axi_master_awuser),      //                                                     .awuser
		.arria10_hps_0_h2f_lw_axi_master_awvalid                    (arria10_hps_0_h2f_lw_axi_master_awvalid),     //                                                     .awvalid
		.arria10_hps_0_h2f_lw_axi_master_awready                    (arria10_hps_0_h2f_lw_axi_master_awready),     //                                                     .awready
		.arria10_hps_0_h2f_lw_axi_master_wid                        (arria10_hps_0_h2f_lw_axi_master_wid),         //                                                     .wid
		.arria10_hps_0_h2f_lw_axi_master_wdata                      (arria10_hps_0_h2f_lw_axi_master_wdata),       //                                                     .wdata
		.arria10_hps_0_h2f_lw_axi_master_wstrb                      (arria10_hps_0_h2f_lw_axi_master_wstrb),       //                                                     .wstrb
		.arria10_hps_0_h2f_lw_axi_master_wlast                      (arria10_hps_0_h2f_lw_axi_master_wlast),       //                                                     .wlast
		.arria10_hps_0_h2f_lw_axi_master_wvalid                     (arria10_hps_0_h2f_lw_axi_master_wvalid),      //                                                     .wvalid
		.arria10_hps_0_h2f_lw_axi_master_wready                     (arria10_hps_0_h2f_lw_axi_master_wready),      //                                                     .wready
		.arria10_hps_0_h2f_lw_axi_master_bid                        (arria10_hps_0_h2f_lw_axi_master_bid),         //                                                     .bid
		.arria10_hps_0_h2f_lw_axi_master_bresp                      (arria10_hps_0_h2f_lw_axi_master_bresp),       //                                                     .bresp
		.arria10_hps_0_h2f_lw_axi_master_bvalid                     (arria10_hps_0_h2f_lw_axi_master_bvalid),      //                                                     .bvalid
		.arria10_hps_0_h2f_lw_axi_master_bready                     (arria10_hps_0_h2f_lw_axi_master_bready),      //                                                     .bready
		.arria10_hps_0_h2f_lw_axi_master_arid                       (arria10_hps_0_h2f_lw_axi_master_arid),        //                                                     .arid
		.arria10_hps_0_h2f_lw_axi_master_araddr                     (arria10_hps_0_h2f_lw_axi_master_araddr),      //                                                     .araddr
		.arria10_hps_0_h2f_lw_axi_master_arlen                      (arria10_hps_0_h2f_lw_axi_master_arlen),       //                                                     .arlen
		.arria10_hps_0_h2f_lw_axi_master_arsize                     (arria10_hps_0_h2f_lw_axi_master_arsize),      //                                                     .arsize
		.arria10_hps_0_h2f_lw_axi_master_arburst                    (arria10_hps_0_h2f_lw_axi_master_arburst),     //                                                     .arburst
		.arria10_hps_0_h2f_lw_axi_master_arlock                     (arria10_hps_0_h2f_lw_axi_master_arlock),      //                                                     .arlock
		.arria10_hps_0_h2f_lw_axi_master_arcache                    (arria10_hps_0_h2f_lw_axi_master_arcache),     //                                                     .arcache
		.arria10_hps_0_h2f_lw_axi_master_arprot                     (arria10_hps_0_h2f_lw_axi_master_arprot),      //                                                     .arprot
		.arria10_hps_0_h2f_lw_axi_master_aruser                     (arria10_hps_0_h2f_lw_axi_master_aruser),      //                                                     .aruser
		.arria10_hps_0_h2f_lw_axi_master_arvalid                    (arria10_hps_0_h2f_lw_axi_master_arvalid),     //                                                     .arvalid
		.arria10_hps_0_h2f_lw_axi_master_arready                    (arria10_hps_0_h2f_lw_axi_master_arready),     //                                                     .arready
		.arria10_hps_0_h2f_lw_axi_master_rid                        (arria10_hps_0_h2f_lw_axi_master_rid),         //                                                     .rid
		.arria10_hps_0_h2f_lw_axi_master_rdata                      (arria10_hps_0_h2f_lw_axi_master_rdata),       //                                                     .rdata
		.arria10_hps_0_h2f_lw_axi_master_rresp                      (arria10_hps_0_h2f_lw_axi_master_rresp),       //                                                     .rresp
		.arria10_hps_0_h2f_lw_axi_master_rlast                      (arria10_hps_0_h2f_lw_axi_master_rlast),       //                                                     .rlast
		.arria10_hps_0_h2f_lw_axi_master_rvalid                     (arria10_hps_0_h2f_lw_axi_master_rvalid),      //                                                     .rvalid
		.arria10_hps_0_h2f_lw_axi_master_rready                     (arria10_hps_0_h2f_lw_axi_master_rready),      //                                                     .rready
		.clk_0_clk_clk                                              (clk_100_clk),                                 //                                            clk_0_clk.clk
		.arria10_hps_0_h2f_lw_axi_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                        // arria10_hps_0_h2f_lw_axi_reset_reset_bridge_in_reset.reset
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset     (hps_fpga_reset_reset),                        //     fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                            (fpga_only_master_master_address),             //                              fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                        (fpga_only_master_master_waitrequest),         //                                                     .waitrequest
		.fpga_only_master_master_byteenable                         (fpga_only_master_master_byteenable),          //                                                     .byteenable
		.fpga_only_master_master_read                               (fpga_only_master_master_read),                //                                                     .read
		.fpga_only_master_master_readdata                           (fpga_only_master_master_readdata),            //                                                     .readdata
		.fpga_only_master_master_readdatavalid                      (fpga_only_master_master_readdatavalid),       //                                                     .readdatavalid
		.fpga_only_master_master_write                              (fpga_only_master_master_write),               //                                                     .write
		.fpga_only_master_master_writedata                          (fpga_only_master_master_writedata),           //                                                     .writedata
		.pb_lwh2f_s0_address                                        (mm_interconnect_1_pb_lwh2f_s0_address),       //                                          pb_lwh2f_s0.address
		.pb_lwh2f_s0_write                                          (mm_interconnect_1_pb_lwh2f_s0_write),         //                                                     .write
		.pb_lwh2f_s0_read                                           (mm_interconnect_1_pb_lwh2f_s0_read),          //                                                     .read
		.pb_lwh2f_s0_readdata                                       (mm_interconnect_1_pb_lwh2f_s0_readdata),      //                                                     .readdata
		.pb_lwh2f_s0_writedata                                      (mm_interconnect_1_pb_lwh2f_s0_writedata),     //                                                     .writedata
		.pb_lwh2f_s0_burstcount                                     (mm_interconnect_1_pb_lwh2f_s0_burstcount),    //                                                     .burstcount
		.pb_lwh2f_s0_byteenable                                     (mm_interconnect_1_pb_lwh2f_s0_byteenable),    //                                                     .byteenable
		.pb_lwh2f_s0_readdatavalid                                  (mm_interconnect_1_pb_lwh2f_s0_readdatavalid), //                                                     .readdatavalid
		.pb_lwh2f_s0_waitrequest                                    (mm_interconnect_1_pb_lwh2f_s0_waitrequest),   //                                                     .waitrequest
		.pb_lwh2f_s0_debugaccess                                    (mm_interconnect_1_pb_lwh2f_s0_debugaccess)    //                                                     .debugaccess
	);

	ghrd_10as066n2_altera_mm_interconnect_161_imhgcbi mm_interconnect_2 (
		.clk_0_clk_clk                              (clk_100_clk),                                           //                            clk_0_clk.clk
		.pb_lwh2f_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                                  // pb_lwh2f_reset_reset_bridge_in_reset.reset
		.pb_lwh2f_m0_address                        (pb_lwh2f_m0_address),                                   //                          pb_lwh2f_m0.address
		.pb_lwh2f_m0_waitrequest                    (pb_lwh2f_m0_waitrequest),                               //                                     .waitrequest
		.pb_lwh2f_m0_burstcount                     (pb_lwh2f_m0_burstcount),                                //                                     .burstcount
		.pb_lwh2f_m0_byteenable                     (pb_lwh2f_m0_byteenable),                                //                                     .byteenable
		.pb_lwh2f_m0_read                           (pb_lwh2f_m0_read),                                      //                                     .read
		.pb_lwh2f_m0_readdata                       (pb_lwh2f_m0_readdata),                                  //                                     .readdata
		.pb_lwh2f_m0_readdatavalid                  (pb_lwh2f_m0_readdatavalid),                             //                                     .readdatavalid
		.pb_lwh2f_m0_write                          (pb_lwh2f_m0_write),                                     //                                     .write
		.pb_lwh2f_m0_writedata                      (pb_lwh2f_m0_writedata),                                 //                                     .writedata
		.pb_lwh2f_m0_debugaccess                    (pb_lwh2f_m0_debugaccess),                               //                                     .debugaccess
		.button_pio_s1_address                      (mm_interconnect_2_button_pio_s1_address),               //                        button_pio_s1.address
		.button_pio_s1_write                        (mm_interconnect_2_button_pio_s1_write),                 //                                     .write
		.button_pio_s1_readdata                     (mm_interconnect_2_button_pio_s1_readdata),              //                                     .readdata
		.button_pio_s1_writedata                    (mm_interconnect_2_button_pio_s1_writedata),             //                                     .writedata
		.button_pio_s1_chipselect                   (mm_interconnect_2_button_pio_s1_chipselect),            //                                     .chipselect
		.dipsw_pio_s1_address                       (mm_interconnect_2_dipsw_pio_s1_address),                //                         dipsw_pio_s1.address
		.dipsw_pio_s1_write                         (mm_interconnect_2_dipsw_pio_s1_write),                  //                                     .write
		.dipsw_pio_s1_readdata                      (mm_interconnect_2_dipsw_pio_s1_readdata),               //                                     .readdata
		.dipsw_pio_s1_writedata                     (mm_interconnect_2_dipsw_pio_s1_writedata),              //                                     .writedata
		.dipsw_pio_s1_chipselect                    (mm_interconnect_2_dipsw_pio_s1_chipselect),             //                                     .chipselect
		.ILC_avalon_slave_address                   (mm_interconnect_2_ilc_avalon_slave_address),            //                     ILC_avalon_slave.address
		.ILC_avalon_slave_write                     (mm_interconnect_2_ilc_avalon_slave_write),              //                                     .write
		.ILC_avalon_slave_read                      (mm_interconnect_2_ilc_avalon_slave_read),               //                                     .read
		.ILC_avalon_slave_readdata                  (mm_interconnect_2_ilc_avalon_slave_readdata),           //                                     .readdata
		.ILC_avalon_slave_writedata                 (mm_interconnect_2_ilc_avalon_slave_writedata),          //                                     .writedata
		.led_pio_s1_address                         (mm_interconnect_2_led_pio_s1_address),                  //                           led_pio_s1.address
		.led_pio_s1_write                           (mm_interconnect_2_led_pio_s1_write),                    //                                     .write
		.led_pio_s1_readdata                        (mm_interconnect_2_led_pio_s1_readdata),                 //                                     .readdata
		.led_pio_s1_writedata                       (mm_interconnect_2_led_pio_s1_writedata),                //                                     .writedata
		.led_pio_s1_chipselect                      (mm_interconnect_2_led_pio_s1_chipselect),               //                                     .chipselect
		.sysid_qsys_0_control_slave_address         (mm_interconnect_2_sysid_qsys_0_control_slave_address),  //           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata        (mm_interconnect_2_sysid_qsys_0_control_slave_readdata)  //                                     .readdata
	);

	ghrd_10as066n2_altera_mm_interconnect_161_kzxwlpi mm_interconnect_3 (
		.arria10_hps_0_f2h_axi_slave_awid                        (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awid),    //                       arria10_hps_0_f2h_axi_slave.awid
		.arria10_hps_0_f2h_axi_slave_awaddr                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awaddr),  //                                                  .awaddr
		.arria10_hps_0_f2h_axi_slave_awlen                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlen),   //                                                  .awlen
		.arria10_hps_0_f2h_axi_slave_awsize                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awsize),  //                                                  .awsize
		.arria10_hps_0_f2h_axi_slave_awburst                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awburst), //                                                  .awburst
		.arria10_hps_0_f2h_axi_slave_awlock                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awlock),  //                                                  .awlock
		.arria10_hps_0_f2h_axi_slave_awcache                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awcache), //                                                  .awcache
		.arria10_hps_0_f2h_axi_slave_awprot                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awprot),  //                                                  .awprot
		.arria10_hps_0_f2h_axi_slave_awuser                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awuser),  //                                                  .awuser
		.arria10_hps_0_f2h_axi_slave_awvalid                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awvalid), //                                                  .awvalid
		.arria10_hps_0_f2h_axi_slave_awready                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_awready), //                                                  .awready
		.arria10_hps_0_f2h_axi_slave_wid                         (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wid),     //                                                  .wid
		.arria10_hps_0_f2h_axi_slave_wdata                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wdata),   //                                                  .wdata
		.arria10_hps_0_f2h_axi_slave_wstrb                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wstrb),   //                                                  .wstrb
		.arria10_hps_0_f2h_axi_slave_wlast                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wlast),   //                                                  .wlast
		.arria10_hps_0_f2h_axi_slave_wvalid                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wvalid),  //                                                  .wvalid
		.arria10_hps_0_f2h_axi_slave_wready                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_wready),  //                                                  .wready
		.arria10_hps_0_f2h_axi_slave_bid                         (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bid),     //                                                  .bid
		.arria10_hps_0_f2h_axi_slave_bresp                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bresp),   //                                                  .bresp
		.arria10_hps_0_f2h_axi_slave_bvalid                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bvalid),  //                                                  .bvalid
		.arria10_hps_0_f2h_axi_slave_bready                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_bready),  //                                                  .bready
		.arria10_hps_0_f2h_axi_slave_arid                        (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arid),    //                                                  .arid
		.arria10_hps_0_f2h_axi_slave_araddr                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_araddr),  //                                                  .araddr
		.arria10_hps_0_f2h_axi_slave_arlen                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlen),   //                                                  .arlen
		.arria10_hps_0_f2h_axi_slave_arsize                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arsize),  //                                                  .arsize
		.arria10_hps_0_f2h_axi_slave_arburst                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arburst), //                                                  .arburst
		.arria10_hps_0_f2h_axi_slave_arlock                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arlock),  //                                                  .arlock
		.arria10_hps_0_f2h_axi_slave_arcache                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arcache), //                                                  .arcache
		.arria10_hps_0_f2h_axi_slave_arprot                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arprot),  //                                                  .arprot
		.arria10_hps_0_f2h_axi_slave_aruser                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_aruser),  //                                                  .aruser
		.arria10_hps_0_f2h_axi_slave_arvalid                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arvalid), //                                                  .arvalid
		.arria10_hps_0_f2h_axi_slave_arready                     (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_arready), //                                                  .arready
		.arria10_hps_0_f2h_axi_slave_rid                         (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rid),     //                                                  .rid
		.arria10_hps_0_f2h_axi_slave_rdata                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rdata),   //                                                  .rdata
		.arria10_hps_0_f2h_axi_slave_rresp                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rresp),   //                                                  .rresp
		.arria10_hps_0_f2h_axi_slave_rlast                       (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rlast),   //                                                  .rlast
		.arria10_hps_0_f2h_axi_slave_rvalid                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rvalid),  //                                                  .rvalid
		.arria10_hps_0_f2h_axi_slave_rready                      (mm_interconnect_3_arria10_hps_0_f2h_axi_slave_rready),  //                                                  .rready
		.clk_0_clk_clk                                           (clk_100_clk),                                           //                                         clk_0_clk.clk
		.arria10_hps_0_f2h_axi_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                                  // arria10_hps_0_f2h_axi_reset_reset_bridge_in_reset.reset
		.hps_only_master_clk_reset_reset_bridge_in_reset_reset   (hps_fpga_reset_reset),                                  //   hps_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_address                          (hps_only_master_master_address),                        //                            hps_only_master_master.address
		.hps_only_master_master_waitrequest                      (hps_only_master_master_waitrequest),                    //                                                  .waitrequest
		.hps_only_master_master_byteenable                       (hps_only_master_master_byteenable),                     //                                                  .byteenable
		.hps_only_master_master_read                             (hps_only_master_master_read),                           //                                                  .read
		.hps_only_master_master_readdata                         (hps_only_master_master_readdata),                       //                                                  .readdata
		.hps_only_master_master_readdatavalid                    (hps_only_master_master_readdatavalid),                  //                                                  .readdatavalid
		.hps_only_master_master_write                            (hps_only_master_master_write),                          //                                                  .write
		.hps_only_master_master_writedata                        (hps_only_master_master_writedata)                       //                                                  .writedata
	);

	ghrd_10as066n2_altera_mm_interconnect_161_srnh6va mm_interconnect_4 (
		.arria10_hps_0_f2sdram0_data_awid                           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awid),    //                          arria10_hps_0_f2sdram0_data.awid
		.arria10_hps_0_f2sdram0_data_awaddr                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awaddr),  //                                                     .awaddr
		.arria10_hps_0_f2sdram0_data_awlen                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlen),   //                                                     .awlen
		.arria10_hps_0_f2sdram0_data_awsize                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awsize),  //                                                     .awsize
		.arria10_hps_0_f2sdram0_data_awburst                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awburst), //                                                     .awburst
		.arria10_hps_0_f2sdram0_data_awlock                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awlock),  //                                                     .awlock
		.arria10_hps_0_f2sdram0_data_awcache                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awcache), //                                                     .awcache
		.arria10_hps_0_f2sdram0_data_awprot                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awprot),  //                                                     .awprot
		.arria10_hps_0_f2sdram0_data_awuser                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awuser),  //                                                     .awuser
		.arria10_hps_0_f2sdram0_data_awvalid                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awvalid), //                                                     .awvalid
		.arria10_hps_0_f2sdram0_data_awready                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_awready), //                                                     .awready
		.arria10_hps_0_f2sdram0_data_wid                            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wid),     //                                                     .wid
		.arria10_hps_0_f2sdram0_data_wdata                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wdata),   //                                                     .wdata
		.arria10_hps_0_f2sdram0_data_wstrb                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wstrb),   //                                                     .wstrb
		.arria10_hps_0_f2sdram0_data_wlast                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wlast),   //                                                     .wlast
		.arria10_hps_0_f2sdram0_data_wvalid                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wvalid),  //                                                     .wvalid
		.arria10_hps_0_f2sdram0_data_wready                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_wready),  //                                                     .wready
		.arria10_hps_0_f2sdram0_data_bid                            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bid),     //                                                     .bid
		.arria10_hps_0_f2sdram0_data_bresp                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bresp),   //                                                     .bresp
		.arria10_hps_0_f2sdram0_data_bvalid                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bvalid),  //                                                     .bvalid
		.arria10_hps_0_f2sdram0_data_bready                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_bready),  //                                                     .bready
		.arria10_hps_0_f2sdram0_data_arid                           (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arid),    //                                                     .arid
		.arria10_hps_0_f2sdram0_data_araddr                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_araddr),  //                                                     .araddr
		.arria10_hps_0_f2sdram0_data_arlen                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlen),   //                                                     .arlen
		.arria10_hps_0_f2sdram0_data_arsize                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arsize),  //                                                     .arsize
		.arria10_hps_0_f2sdram0_data_arburst                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arburst), //                                                     .arburst
		.arria10_hps_0_f2sdram0_data_arlock                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arlock),  //                                                     .arlock
		.arria10_hps_0_f2sdram0_data_arcache                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arcache), //                                                     .arcache
		.arria10_hps_0_f2sdram0_data_arprot                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arprot),  //                                                     .arprot
		.arria10_hps_0_f2sdram0_data_aruser                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_aruser),  //                                                     .aruser
		.arria10_hps_0_f2sdram0_data_arvalid                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arvalid), //                                                     .arvalid
		.arria10_hps_0_f2sdram0_data_arready                        (mm_interconnect_4_arria10_hps_0_f2sdram0_data_arready), //                                                     .arready
		.arria10_hps_0_f2sdram0_data_rid                            (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rid),     //                                                     .rid
		.arria10_hps_0_f2sdram0_data_rdata                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rdata),   //                                                     .rdata
		.arria10_hps_0_f2sdram0_data_rresp                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rresp),   //                                                     .rresp
		.arria10_hps_0_f2sdram0_data_rlast                          (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rlast),   //                                                     .rlast
		.arria10_hps_0_f2sdram0_data_rvalid                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rvalid),  //                                                     .rvalid
		.arria10_hps_0_f2sdram0_data_rready                         (mm_interconnect_4_arria10_hps_0_f2sdram0_data_rready),  //                                                     .rready
		.clk_0_clk_clk                                              (clk_100_clk),                                           //                                            clk_0_clk.clk
		.arria10_hps_0_f2sdram0_reset_reset_bridge_in_reset_reset   (hps_fpga_reset_reset),                                  //   arria10_hps_0_f2sdram0_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master1_clk_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                                  // f2sdram_only_master1_clk_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master1_master_address                        (f2sdram_only_master1_master_address),                   //                          f2sdram_only_master1_master.address
		.f2sdram_only_master1_master_waitrequest                    (f2sdram_only_master1_master_waitrequest),               //                                                     .waitrequest
		.f2sdram_only_master1_master_byteenable                     (f2sdram_only_master1_master_byteenable),                //                                                     .byteenable
		.f2sdram_only_master1_master_read                           (f2sdram_only_master1_master_read),                      //                                                     .read
		.f2sdram_only_master1_master_readdata                       (f2sdram_only_master1_master_readdata),                  //                                                     .readdata
		.f2sdram_only_master1_master_readdatavalid                  (f2sdram_only_master1_master_readdatavalid),             //                                                     .readdatavalid
		.f2sdram_only_master1_master_write                          (f2sdram_only_master1_master_write),                     //                                                     .write
		.f2sdram_only_master1_master_writedata                      (f2sdram_only_master1_master_writedata)                  //                                                     .writedata
	);

	ghrd_10as066n2_altera_mm_interconnect_161_a4dxs3y mm_interconnect_5 (
		.arria10_hps_0_f2sdram2_data_awid                          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awid),    //                         arria10_hps_0_f2sdram2_data.awid
		.arria10_hps_0_f2sdram2_data_awaddr                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awaddr),  //                                                    .awaddr
		.arria10_hps_0_f2sdram2_data_awlen                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlen),   //                                                    .awlen
		.arria10_hps_0_f2sdram2_data_awsize                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awsize),  //                                                    .awsize
		.arria10_hps_0_f2sdram2_data_awburst                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awburst), //                                                    .awburst
		.arria10_hps_0_f2sdram2_data_awlock                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awlock),  //                                                    .awlock
		.arria10_hps_0_f2sdram2_data_awcache                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awcache), //                                                    .awcache
		.arria10_hps_0_f2sdram2_data_awprot                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awprot),  //                                                    .awprot
		.arria10_hps_0_f2sdram2_data_awuser                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awuser),  //                                                    .awuser
		.arria10_hps_0_f2sdram2_data_awvalid                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awvalid), //                                                    .awvalid
		.arria10_hps_0_f2sdram2_data_awready                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_awready), //                                                    .awready
		.arria10_hps_0_f2sdram2_data_wid                           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wid),     //                                                    .wid
		.arria10_hps_0_f2sdram2_data_wdata                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wdata),   //                                                    .wdata
		.arria10_hps_0_f2sdram2_data_wstrb                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wstrb),   //                                                    .wstrb
		.arria10_hps_0_f2sdram2_data_wlast                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wlast),   //                                                    .wlast
		.arria10_hps_0_f2sdram2_data_wvalid                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wvalid),  //                                                    .wvalid
		.arria10_hps_0_f2sdram2_data_wready                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_wready),  //                                                    .wready
		.arria10_hps_0_f2sdram2_data_bid                           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bid),     //                                                    .bid
		.arria10_hps_0_f2sdram2_data_bresp                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bresp),   //                                                    .bresp
		.arria10_hps_0_f2sdram2_data_bvalid                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bvalid),  //                                                    .bvalid
		.arria10_hps_0_f2sdram2_data_bready                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_bready),  //                                                    .bready
		.arria10_hps_0_f2sdram2_data_arid                          (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arid),    //                                                    .arid
		.arria10_hps_0_f2sdram2_data_araddr                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_araddr),  //                                                    .araddr
		.arria10_hps_0_f2sdram2_data_arlen                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlen),   //                                                    .arlen
		.arria10_hps_0_f2sdram2_data_arsize                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arsize),  //                                                    .arsize
		.arria10_hps_0_f2sdram2_data_arburst                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arburst), //                                                    .arburst
		.arria10_hps_0_f2sdram2_data_arlock                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arlock),  //                                                    .arlock
		.arria10_hps_0_f2sdram2_data_arcache                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arcache), //                                                    .arcache
		.arria10_hps_0_f2sdram2_data_arprot                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arprot),  //                                                    .arprot
		.arria10_hps_0_f2sdram2_data_aruser                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_aruser),  //                                                    .aruser
		.arria10_hps_0_f2sdram2_data_arvalid                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arvalid), //                                                    .arvalid
		.arria10_hps_0_f2sdram2_data_arready                       (mm_interconnect_5_arria10_hps_0_f2sdram2_data_arready), //                                                    .arready
		.arria10_hps_0_f2sdram2_data_rid                           (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rid),     //                                                    .rid
		.arria10_hps_0_f2sdram2_data_rdata                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rdata),   //                                                    .rdata
		.arria10_hps_0_f2sdram2_data_rresp                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rresp),   //                                                    .rresp
		.arria10_hps_0_f2sdram2_data_rlast                         (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rlast),   //                                                    .rlast
		.arria10_hps_0_f2sdram2_data_rvalid                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rvalid),  //                                                    .rvalid
		.arria10_hps_0_f2sdram2_data_rready                        (mm_interconnect_5_arria10_hps_0_f2sdram2_data_rready),  //                                                    .rready
		.clk_0_clk_clk                                             (clk_100_clk),                                           //                                           clk_0_clk.clk
		.arria10_hps_0_f2sdram2_reset_reset_bridge_in_reset_reset  (hps_fpga_reset_reset),                                  //  arria10_hps_0_f2sdram2_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset (hps_fpga_reset_reset),                                  // f2sdram_only_master_clk_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_address                        (f2sdram_only_master_master_address),                    //                          f2sdram_only_master_master.address
		.f2sdram_only_master_master_waitrequest                    (f2sdram_only_master_master_waitrequest),                //                                                    .waitrequest
		.f2sdram_only_master_master_byteenable                     (f2sdram_only_master_master_byteenable),                 //                                                    .byteenable
		.f2sdram_only_master_master_read                           (f2sdram_only_master_master_read),                       //                                                    .read
		.f2sdram_only_master_master_readdata                       (f2sdram_only_master_master_readdata),                   //                                                    .readdata
		.f2sdram_only_master_master_readdatavalid                  (f2sdram_only_master_master_readdatavalid),              //                                                    .readdatavalid
		.f2sdram_only_master_master_write                          (f2sdram_only_master_master_write),                      //                                                    .write
		.f2sdram_only_master_master_writedata                      (f2sdram_only_master_master_writedata)                   //                                                    .writedata
	);

	ghrd_10as066n2_altera_irq_mapper_161_nvquryy irq_mapper (
		.clk           (clk_100_clk),              //       clk.clk
		.reset         (hps_fpga_reset_reset),     // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (ilc_irq_irq)               //    sender.irq
	);

	ghrd_10as066n2_altera_irq_mapper_161_43ijldi irq_mapper_001 (
		.clk           (),                           //       clk.clk
		.reset         (),                           // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),   // receiver1.irq
		.sender_irq    (arria10_hps_0_f2h_irq0_irq)  //    sender.irq
	);

	ghrd_10as066n2_altera_irq_mapper_161_kbptgda irq_mapper_002 (
		.clk        (),                           //       clk.clk
		.reset      (),                           // clk_reset.reset
		.sender_irq (arria10_hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~arria10_hps_0_h2f_reset_reset),     // reset_in1.reset
		.clk            (clk_100_clk),                        //       clk.clk
		.reset_out      (hps_fpga_reset_reset),               // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~arria10_hps_0_h2f_reset_reset),     // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~arria10_hps_0_h2f_reset_reset),     // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~arria10_hps_0_h2f_reset_reset),     // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~arria10_hps_0_h2f_reset_reset),     // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
