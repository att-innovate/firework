// extender_8to32.v

module extender_8to32 (
		// TODO: define ports
	);
	
	// TODO: define extender logic
	
endmodule
