// extender_8to32.v

module extender_8to32 (
		// clock, reset inputs
		input  wire        clk,
		input  wire        reset

		// TODO: define ports
	);
	
	// TODO: define extender logic
	
endmodule
