// raw_data_out_index.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module raw_data_out_index (
		input  wire [9:0] data,  //  fifo_input.datain
		input  wire       wrreq, //            .wrreq
		input  wire       rdreq, //            .rdreq
		input  wire       clock, //            .clk
		input  wire       sclr,  //            .sclr
		output wire [9:0] q      // fifo_output.dataout
	);

	raw_data_out_index_fifo_171_z22fama fifo_0 (
		.data  (data),  //  fifo_input.datain
		.wrreq (wrreq), //            .wrreq
		.rdreq (rdreq), //            .rdreq
		.clock (clock), //            .clk
		.sclr  (sclr),  //            .sclr
		.q     (q)      // fifo_output.dataout
	);

endmodule
