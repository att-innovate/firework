
module varint_in_size (
	data,
	wrreq,
	rdreq,
	clock,
	sclr,
	q);	

	input		data;
	input		wrreq;
	input		rdreq;
	input		clock;
	input		sclr;
	output		q;
endmodule
