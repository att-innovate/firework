// varint_in_size.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module varint_in_size (
		input  wire  data,  //  fifo_input.datain
		input  wire  wrreq, //            .wrreq
		input  wire  rdreq, //            .rdreq
		input  wire  clock, //            .clk
		input  wire  sclr,  //            .sclr
		output wire  q      // fifo_output.dataout
	);

	varint_in_size_fifo_160_sjmeklq fifo_0 (
		.data  (data),  //  fifo_input.datain
		.wrreq (wrreq), //            .wrreq
		.rdreq (rdreq), //            .rdreq
		.clock (clock), //            .clk
		.sclr  (sclr),  //            .sclr
		.q     (q)      // fifo_output.dataout
	);

endmodule
