module varint_encoder_top (
	input wire [31:0]	data,
	input wire			valid,
	output wire			ready
);


endmodule
