// in_fifo.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module in_fifo (
		input  wire [31:0] data,  //  fifo_input.datain
		input  wire        wrreq, //            .wrreq
		input  wire        rdreq, //            .rdreq
		input  wire        clock, //            .clk
		input  wire        sclr,  //            .sclr
		output wire [31:0] q,     // fifo_output.dataout
		output wire [9:0]  usedw, //            .usedw
		output wire        full,  //            .full
		output wire        empty  //            .empty
	);

	in_fifo_fifo_160_mnfmh2i fifo_0 (
		.data  (data),  //  fifo_input.datain
		.wrreq (wrreq), //            .wrreq
		.rdreq (rdreq), //            .rdreq
		.clock (clock), //            .clk
		.sclr  (sclr),  //            .sclr
		.q     (q),     // fifo_output.dataout
		.usedw (usedw), //            .usedw
		.full  (full),  //            .full
		.empty (empty)  //            .empty
	);

endmodule
